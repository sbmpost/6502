module MEMORY(
  input CLK,
  input WE,
  input[15:0] Address,
  input[7:0] DataIn,
  output reg[7:0] DataOut
);

//  reg [7:0] s_mem_contents[65535:0];
  reg [7:0] s_mem_contents[16383:0];
  parameter b_lo = 8'h00;
  parameter b_hi = 8'h04;
  parameter base = {b_hi, b_lo};

  initial begin

`ifdef VERILATOR

      // LDX #07 (x=7)
      s_mem_contents[base + 00] = 8'ha2;
      s_mem_contents[base + 01] = 8'h07;
      // LDY #08 (y=8)
      s_mem_contents[base + 02] = 8'ha0;
      s_mem_contents[base + 03] = 8'h08;
      // LDA $00ff,y (y=8)
      s_mem_contents[base + 04] = 8'hb9;
      s_mem_contents[base + 05] = 8'hff;
      s_mem_contents[base + 06] = 8'h00;
      // LDA $0108,y (y=8)
      s_mem_contents[base + 07] = 8'hb9;
      s_mem_contents[base + 08] = 8'h08;
      s_mem_contents[base + 09] = 8'h01;
      // LDA $01f0,x (x=7)
      s_mem_contents[base + 10] = 8'hbd;
      s_mem_contents[base + 11] = 8'hf0;
      s_mem_contents[base + 12] = 8'h01;
      // LDA $30,x (x=7)
      s_mem_contents[base + 13] = 8'hb5;
      s_mem_contents[base + 14] = 8'h30;
      // LDA $40,x (x=7)
      s_mem_contents[base + 15] = 8'hb5;
      s_mem_contents[base + 16] = 8'h40;
      // LDA $ff,x (x=7), should access $0006
      s_mem_contents[base + 17] = 8'hb5;
      s_mem_contents[base + 18] = 8'hff;
      // LDA $0110
      s_mem_contents[base + 19] = 8'had;
      s_mem_contents[base + 20] = 8'h10;
      s_mem_contents[base + 21] = 8'h01;
      // LDA $37
      s_mem_contents[base + 22] = 8'ha5;
      s_mem_contents[base + 23] = 8'h37;
      // LDA ($1e),y (y=8, $1e=fc, $1f=02), should access $0304
      s_mem_contents[base + 24] = 8'hb1;
      s_mem_contents[base + 25] = 8'h1e;
      // JMP $0021
      s_mem_contents[base + 26] = 8'h4c;
      s_mem_contents[base + 27] = 8'h21;
      s_mem_contents[base + 28] = b_hi;

      // data
      s_mem_contents[11] = 8'hf0;
      s_mem_contents[25] = 8'h1e;
      s_mem_contents[29] = 8'h00;
      s_mem_contents[30] = 8'hfc;
      s_mem_contents[31] = 8'h02;
      s_mem_contents[32] = 8'hfe;

      // STA $0108,y (y=8)
      s_mem_contents[base + 33] = 8'h99;
      s_mem_contents[base + 34] = 8'h08;
      s_mem_contents[base + 35] = 8'h01;
      // LDA #19
      s_mem_contents[base + 36] = 8'ha9;
      s_mem_contents[base + 37] = 8'h19;
      // LDA $0108,y (y=8)
      s_mem_contents[base + 38] = 8'hb9;
      s_mem_contents[base + 39] = 8'h08;
      s_mem_contents[base + 40] = 8'h01;
      // LDA #20
      s_mem_contents[base + 41] = 8'ha9;
      s_mem_contents[base + 42] = 8'h20;
      // STA $00ff,x (x=7) $0106
      s_mem_contents[base + 43] = 8'h9d;
      s_mem_contents[base + 44] = 8'hff;
      s_mem_contents[base + 45] = 8'h00;
      // LDA #21
      s_mem_contents[base + 46] = 8'ha9;
      s_mem_contents[base + 47] = 8'h21;
      // LDA $00ff,x (x=7) $0106
      s_mem_contents[base + 48] = 8'hbd;
      s_mem_contents[base + 49] = 8'hff;
      s_mem_contents[base + 50] = 8'h00;
      // JMP $0305
      s_mem_contents[base + 51] = 8'h4c;
      s_mem_contents[base + 52] = 8'h05;
      s_mem_contents[base + 53] = 8'h03+b_hi;

      // data
      s_mem_contents[55] = 8'hdd;
      s_mem_contents[71] = 8'hee;
      s_mem_contents[263] = 8'haa;
      s_mem_contents[272] = 8'hbb;
      s_mem_contents[503] = 8'hcc;
      s_mem_contents[512] = 8'h03+b_hi;

      // LDX $01ab,y
      s_mem_contents[base + 724] = 8'hbe; // $02d4
      s_mem_contents[base + 725] = 8'hab;
      s_mem_contents[base + 726] = 8'h01;
      // STX $77,y
      s_mem_contents[base + 727] = 8'h96;
      s_mem_contents[base + 728] = 8'h77;
      // DEX
      s_mem_contents[base + 729] = 8'hca;
      // LDA ($20,x)
      s_mem_contents[base + 730] = 8'ha1;
      s_mem_contents[base + 731] = 8'h20;
      // BVC $74
      s_mem_contents[base + 732] = 8'h50;
      s_mem_contents[base + 733] = 8'h74; // $02dc

      // data
      s_mem_contents[766] = 8'h33; // $02fe
      s_mem_contents[767] = 8'h10; // $02ff
      s_mem_contents[772] = 8'hff; // $0304
      s_mem_contents[773] = 8'he8; // $0305

      // INX
      s_mem_contents[base + 773] = 8'he8;
      // INY
      s_mem_contents[base + 774] = 8'hc8;
      // DEX
      s_mem_contents[base + 775] = 8'hca;
      // DEY
      s_mem_contents[base + 776] = 8'h88;
      // JMP ($02ff)
      s_mem_contents[base + 777] = 8'h6c;
      s_mem_contents[base + 778] = 8'hff;
      s_mem_contents[base + 779] = 8'h02;
      s_mem_contents[base + 780] = 8'h00;
      s_mem_contents[base + 781] = 8'h00;
      s_mem_contents[base + 782] = 8'h00;
      s_mem_contents[base + 783] = 8'h00;
      // TXA
      s_mem_contents[base + 784] = 8'h8a;
      // TYA
      s_mem_contents[base + 785] = 8'h98;
      // TAX
      s_mem_contents[base + 786] = 8'haa;
      // INY
      s_mem_contents[base + 787] = 8'hc8;
      // TAY
      s_mem_contents[base + 788] = 8'ha8;
      // INY
      s_mem_contents[base + 789] = 8'hc8;
      // ORA $02f7,x (x=8)
      s_mem_contents[base + 790] = 8'h1d;
      s_mem_contents[base + 791] = 8'hf7;
      s_mem_contents[base + 792] = 8'h02;
      // AND $0b
      s_mem_contents[base + 793] = 8'h25;
      s_mem_contents[base + 794] = 8'h0b;
      // EOR ($1e),y (y=8)
      s_mem_contents[base + 795] = 8'h51;
      s_mem_contents[base + 796] = 8'h1e;
      // ADC #08
      s_mem_contents[base + 797] = 8'h69;
      s_mem_contents[base + 798] = 8'h08;
      // ADC $02fc,x (x=8)
      s_mem_contents[base + 799] = 8'h7d;
      s_mem_contents[base + 800] = 8'hfc;
      s_mem_contents[base + 801] = 8'h02;
      // SBC #44
      s_mem_contents[base + 802] = 8'he9;
      s_mem_contents[base + 803] = 8'h44;
      // CPY $01
      s_mem_contents[base + 804] = 8'hc4;
      s_mem_contents[base + 805] = 8'h01;
      // CPX $0304
      s_mem_contents[base + 806] = 8'hec;
      s_mem_contents[base + 807] = 8'h04;
      s_mem_contents[base + 808] = 8'h03;
      // CMP ($1e),y
      s_mem_contents[base + 809] = 8'hd1;
      s_mem_contents[base + 810] = 8'h1e;
      // INC $02ff
      s_mem_contents[base + 811] = 8'hee;
      s_mem_contents[base + 812] = 8'hff;
      s_mem_contents[base + 813] = 8'h02;
      // LDX $02ff
      s_mem_contents[base + 814] = 8'hae;
      s_mem_contents[base + 815] = 8'hff;
      s_mem_contents[base + 816] = 8'h02;
      // DEC $08,x
      s_mem_contents[base + 817] = 8'hd6;
      s_mem_contents[base + 818] = 8'h08;
      // LDA #81
      s_mem_contents[base + 819] = 8'ha9;
      s_mem_contents[base + 820] = 8'h81;
      // LSR A
      s_mem_contents[base + 821] = 8'h4a;
      // ROL A
      s_mem_contents[base + 822] = 8'h2a;
      // ASL A
      s_mem_contents[base + 823] = 8'h0a;
      // ROR A
      s_mem_contents[base + 824] = 8'h6a;
      // LDY $08,x
      s_mem_contents[base + 825] = 8'hb4;
      s_mem_contents[base + 826] = 8'h08;
      // LSR $08,x
      s_mem_contents[base + 827] = 8'h56;
      s_mem_contents[base + 828] = 8'h08;
      // LDY $08,x
      s_mem_contents[base + 829] = 8'hb4;
      s_mem_contents[base + 830] = 8'h08;
      // ASL $08,x
      s_mem_contents[base + 831] = 8'h16;
      s_mem_contents[base + 832] = 8'h08;
      // LDY $08,x
      s_mem_contents[base + 833] = 8'hb4;
      s_mem_contents[base + 834] = 8'h08;
      // ROR $08,x
      s_mem_contents[base + 835] = 8'h76;
      s_mem_contents[base + 836] = 8'h08;
      // LDY $08,x
      s_mem_contents[base + 837] = 8'hb4;
      s_mem_contents[base + 838] = 8'h08;
      // ROL $08,x
      s_mem_contents[base + 839] = 8'h36;
      s_mem_contents[base + 840] = 8'h08;
      // LDY $08,x
      s_mem_contents[base + 841] = 8'hb4;
      s_mem_contents[base + 842] = 8'h08;
      // SEC
      s_mem_contents[base + 843] = 8'h38;
      // CLC
      s_mem_contents[base + 844] = 8'h18;
      // CLV
      s_mem_contents[base + 845] = 8'hb8;
      // BVS $02
      s_mem_contents[base + 846] = 8'h70; // $034e
      s_mem_contents[base + 847] = 8'h02; // $034f
      // BVC $80
      s_mem_contents[base + 848] = 8'h50; // $0350
      s_mem_contents[base + 849] = 8'h80; // $0351
      // INX
      s_mem_contents[base + 850] = 8'he8;
      // DEX
      s_mem_contents[base + 851] = 8'hca;
      // LDA #01
      s_mem_contents[base + 852] = 8'ha9;
      s_mem_contents[base + 853] = 8'h01;
      // TXA
      s_mem_contents[base + 854] = 8'h8a;
      // TSX
      s_mem_contents[base + 855] = 8'hba;
      // NOP
      s_mem_contents[base + 856] = 8'hea;
      // PHP
      s_mem_contents[base + 857] = 8'h08;
      // PHA
      s_mem_contents[base + 858] = 8'h48;
      // PLP
      s_mem_contents[base + 859] = 8'h28;
      // PLA
      s_mem_contents[base + 860] = 8'h68;
      // NOP
      s_mem_contents[base + 861] = 8'hea;
      // JSR $0364
      s_mem_contents[base + 862] = 8'h20; // $035e
      s_mem_contents[base + 863] = 8'h64; // $035f
      s_mem_contents[base + 864] = 8'h03+b_hi; // $0360
      // JMP $0366
      s_mem_contents[base + 865] = 8'h4c; // $0361
      s_mem_contents[base + 866] = 8'h66; // $0362
      s_mem_contents[base + 867] = 8'h03+b_hi; // $0363
      // NOP
      s_mem_contents[base + 868] = 8'hea; // $0364
      // RTS
      s_mem_contents[base + 869] = 8'h60; // $0365
      // NOP
      s_mem_contents[base + 870] = 8'hea; // $0366

`else

s_mem_contents[14'h0000] = 8'h00;
s_mem_contents[14'h0001] = 8'h00;
s_mem_contents[14'h0002] = 8'h00;
s_mem_contents[14'h0003] = 8'h00;
s_mem_contents[14'h0004] = 8'h00;
s_mem_contents[14'h0005] = 8'h00;
s_mem_contents[14'h0006] = 8'h00;
s_mem_contents[14'h0007] = 8'h00;
s_mem_contents[14'h0008] = 8'h00;
s_mem_contents[14'h0009] = 8'hc3;
s_mem_contents[14'h000a] = 8'h82;
s_mem_contents[14'h000b] = 8'h41;
s_mem_contents[14'h000c] = 8'h00;
s_mem_contents[14'h000d] = 8'h7f;
s_mem_contents[14'h000e] = 8'h00;
s_mem_contents[14'h000f] = 8'h1f;
s_mem_contents[14'h0010] = 8'h71;
s_mem_contents[14'h0011] = 8'h80;
s_mem_contents[14'h0012] = 8'h0f;
s_mem_contents[14'h0013] = 8'hff;
s_mem_contents[14'h0014] = 8'h7f;
s_mem_contents[14'h0015] = 8'h80;
s_mem_contents[14'h0016] = 8'hff;
s_mem_contents[14'h0017] = 8'h0f;
s_mem_contents[14'h0018] = 8'h8f;
s_mem_contents[14'h0019] = 8'h8f;
s_mem_contents[14'h001a] = 8'h17;
s_mem_contents[14'h001b] = 8'h02;
s_mem_contents[14'h001c] = 8'h18;
s_mem_contents[14'h001d] = 8'h02;
s_mem_contents[14'h001e] = 8'h19;
s_mem_contents[14'h001f] = 8'h02;
s_mem_contents[14'h0020] = 8'h1a;
s_mem_contents[14'h0021] = 8'h02;
s_mem_contents[14'h0022] = 8'h1b;
s_mem_contents[14'h0023] = 8'h02;
s_mem_contents[14'h0024] = 8'h1f;
s_mem_contents[14'h0025] = 8'h01;
s_mem_contents[14'h0026] = 8'h03;
s_mem_contents[14'h0027] = 8'h02;
s_mem_contents[14'h0028] = 8'h04;
s_mem_contents[14'h0029] = 8'h02;
s_mem_contents[14'h002a] = 8'h05;
s_mem_contents[14'h002b] = 8'h02;
s_mem_contents[14'h002c] = 8'h06;
s_mem_contents[14'h002d] = 8'h02;
s_mem_contents[14'h002e] = 8'h0b;
s_mem_contents[14'h002f] = 8'h01;
s_mem_contents[14'h0030] = 8'h4e;
s_mem_contents[14'h0031] = 8'h02;
s_mem_contents[14'h0032] = 8'h4f;
s_mem_contents[14'h0033] = 8'h02;
s_mem_contents[14'h0034] = 8'h50;
s_mem_contents[14'h0035] = 8'h02;
s_mem_contents[14'h0036] = 8'h51;
s_mem_contents[14'h0037] = 8'h02;
s_mem_contents[14'h0038] = 8'h52;
s_mem_contents[14'h0039] = 8'h02;
s_mem_contents[14'h003a] = 8'h53;
s_mem_contents[14'h003b] = 8'h02;
s_mem_contents[14'h003c] = 8'h54;
s_mem_contents[14'h003d] = 8'h02;
s_mem_contents[14'h003e] = 8'h55;
s_mem_contents[14'h003f] = 8'h02;
s_mem_contents[14'h0040] = 8'h4a;
s_mem_contents[14'h0041] = 8'h02;
s_mem_contents[14'h0042] = 8'h4b;
s_mem_contents[14'h0043] = 8'h02;
s_mem_contents[14'h0044] = 8'h4c;
s_mem_contents[14'h0045] = 8'h02;
s_mem_contents[14'h0046] = 8'h4d;
s_mem_contents[14'h0047] = 8'h02;
s_mem_contents[14'h0048] = 8'h03;
s_mem_contents[14'h0049] = 8'h02;
s_mem_contents[14'h004a] = 8'h04;
s_mem_contents[14'h004b] = 8'h02;
s_mem_contents[14'h004c] = 8'h04;
s_mem_contents[14'h004d] = 8'h01;
s_mem_contents[14'h004e] = 8'h05;
s_mem_contents[14'h004f] = 8'h01;
s_mem_contents[14'h0050] = 8'hff;
s_mem_contents[14'h0051] = 8'hff;
s_mem_contents[14'h0052] = 8'hff;
s_mem_contents[14'h0053] = 8'hff;
s_mem_contents[14'h0054] = 8'hff;
s_mem_contents[14'h0055] = 8'hff;
s_mem_contents[14'h0056] = 8'hff;
s_mem_contents[14'h0057] = 8'hff;
s_mem_contents[14'h0058] = 8'hff;
s_mem_contents[14'h0059] = 8'hff;
s_mem_contents[14'h005a] = 8'hff;
s_mem_contents[14'h005b] = 8'hff;
s_mem_contents[14'h005c] = 8'hff;
s_mem_contents[14'h005d] = 8'hff;
s_mem_contents[14'h005e] = 8'hff;
s_mem_contents[14'h005f] = 8'hff;
s_mem_contents[14'h0060] = 8'hff;
s_mem_contents[14'h0061] = 8'hff;
s_mem_contents[14'h0062] = 8'hff;
s_mem_contents[14'h0063] = 8'hff;
s_mem_contents[14'h0064] = 8'hff;
s_mem_contents[14'h0065] = 8'hff;
s_mem_contents[14'h0066] = 8'hff;
s_mem_contents[14'h0067] = 8'hff;
s_mem_contents[14'h0068] = 8'hff;
s_mem_contents[14'h0069] = 8'hff;
s_mem_contents[14'h006a] = 8'hff;
s_mem_contents[14'h006b] = 8'hff;
s_mem_contents[14'h006c] = 8'hff;
s_mem_contents[14'h006d] = 8'hff;
s_mem_contents[14'h006e] = 8'hff;
s_mem_contents[14'h006f] = 8'hff;
s_mem_contents[14'h0070] = 8'hff;
s_mem_contents[14'h0071] = 8'hff;
s_mem_contents[14'h0072] = 8'hff;
s_mem_contents[14'h0073] = 8'hff;
s_mem_contents[14'h0074] = 8'hff;
s_mem_contents[14'h0075] = 8'hff;
s_mem_contents[14'h0076] = 8'hff;
s_mem_contents[14'h0077] = 8'hff;
s_mem_contents[14'h0078] = 8'hff;
s_mem_contents[14'h0079] = 8'hff;
s_mem_contents[14'h007a] = 8'hff;
s_mem_contents[14'h007b] = 8'hff;
s_mem_contents[14'h007c] = 8'hff;
s_mem_contents[14'h007d] = 8'hff;
s_mem_contents[14'h007e] = 8'hff;
s_mem_contents[14'h007f] = 8'hff;
s_mem_contents[14'h0080] = 8'hff;
s_mem_contents[14'h0081] = 8'hff;
s_mem_contents[14'h0082] = 8'hff;
s_mem_contents[14'h0083] = 8'hff;
s_mem_contents[14'h0084] = 8'hff;
s_mem_contents[14'h0085] = 8'hff;
s_mem_contents[14'h0086] = 8'hff;
s_mem_contents[14'h0087] = 8'hff;
s_mem_contents[14'h0088] = 8'hff;
s_mem_contents[14'h0089] = 8'hff;
s_mem_contents[14'h008a] = 8'hff;
s_mem_contents[14'h008b] = 8'hff;
s_mem_contents[14'h008c] = 8'hff;
s_mem_contents[14'h008d] = 8'hff;
s_mem_contents[14'h008e] = 8'hff;
s_mem_contents[14'h008f] = 8'hff;
s_mem_contents[14'h0090] = 8'hff;
s_mem_contents[14'h0091] = 8'hff;
s_mem_contents[14'h0092] = 8'hff;
s_mem_contents[14'h0093] = 8'hff;
s_mem_contents[14'h0094] = 8'hff;
s_mem_contents[14'h0095] = 8'hff;
s_mem_contents[14'h0096] = 8'hff;
s_mem_contents[14'h0097] = 8'hff;
s_mem_contents[14'h0098] = 8'hff;
s_mem_contents[14'h0099] = 8'hff;
s_mem_contents[14'h009a] = 8'hff;
s_mem_contents[14'h009b] = 8'hff;
s_mem_contents[14'h009c] = 8'hff;
s_mem_contents[14'h009d] = 8'hff;
s_mem_contents[14'h009e] = 8'hff;
s_mem_contents[14'h009f] = 8'hff;
s_mem_contents[14'h00a0] = 8'hff;
s_mem_contents[14'h00a1] = 8'hff;
s_mem_contents[14'h00a2] = 8'hff;
s_mem_contents[14'h00a3] = 8'hff;
s_mem_contents[14'h00a4] = 8'hff;
s_mem_contents[14'h00a5] = 8'hff;
s_mem_contents[14'h00a6] = 8'hff;
s_mem_contents[14'h00a7] = 8'hff;
s_mem_contents[14'h00a8] = 8'hff;
s_mem_contents[14'h00a9] = 8'hff;
s_mem_contents[14'h00aa] = 8'hff;
s_mem_contents[14'h00ab] = 8'hff;
s_mem_contents[14'h00ac] = 8'hff;
s_mem_contents[14'h00ad] = 8'hff;
s_mem_contents[14'h00ae] = 8'hff;
s_mem_contents[14'h00af] = 8'hff;
s_mem_contents[14'h00b0] = 8'hff;
s_mem_contents[14'h00b1] = 8'hff;
s_mem_contents[14'h00b2] = 8'hff;
s_mem_contents[14'h00b3] = 8'hff;
s_mem_contents[14'h00b4] = 8'hff;
s_mem_contents[14'h00b5] = 8'hff;
s_mem_contents[14'h00b6] = 8'hff;
s_mem_contents[14'h00b7] = 8'hff;
s_mem_contents[14'h00b8] = 8'hff;
s_mem_contents[14'h00b9] = 8'hff;
s_mem_contents[14'h00ba] = 8'hff;
s_mem_contents[14'h00bb] = 8'hff;
s_mem_contents[14'h00bc] = 8'hff;
s_mem_contents[14'h00bd] = 8'hff;
s_mem_contents[14'h00be] = 8'hff;
s_mem_contents[14'h00bf] = 8'hff;
s_mem_contents[14'h00c0] = 8'hff;
s_mem_contents[14'h00c1] = 8'hff;
s_mem_contents[14'h00c2] = 8'hff;
s_mem_contents[14'h00c3] = 8'hff;
s_mem_contents[14'h00c4] = 8'hff;
s_mem_contents[14'h00c5] = 8'hff;
s_mem_contents[14'h00c6] = 8'hff;
s_mem_contents[14'h00c7] = 8'hff;
s_mem_contents[14'h00c8] = 8'hff;
s_mem_contents[14'h00c9] = 8'hff;
s_mem_contents[14'h00ca] = 8'hff;
s_mem_contents[14'h00cb] = 8'hff;
s_mem_contents[14'h00cc] = 8'hff;
s_mem_contents[14'h00cd] = 8'hff;
s_mem_contents[14'h00ce] = 8'hff;
s_mem_contents[14'h00cf] = 8'hff;
s_mem_contents[14'h00d0] = 8'hff;
s_mem_contents[14'h00d1] = 8'hff;
s_mem_contents[14'h00d2] = 8'hff;
s_mem_contents[14'h00d3] = 8'hff;
s_mem_contents[14'h00d4] = 8'hff;
s_mem_contents[14'h00d5] = 8'hff;
s_mem_contents[14'h00d6] = 8'hff;
s_mem_contents[14'h00d7] = 8'hff;
s_mem_contents[14'h00d8] = 8'hff;
s_mem_contents[14'h00d9] = 8'hff;
s_mem_contents[14'h00da] = 8'hff;
s_mem_contents[14'h00db] = 8'hff;
s_mem_contents[14'h00dc] = 8'hff;
s_mem_contents[14'h00dd] = 8'hff;
s_mem_contents[14'h00de] = 8'hff;
s_mem_contents[14'h00df] = 8'hff;
s_mem_contents[14'h00e0] = 8'hff;
s_mem_contents[14'h00e1] = 8'hff;
s_mem_contents[14'h00e2] = 8'hff;
s_mem_contents[14'h00e3] = 8'hff;
s_mem_contents[14'h00e4] = 8'hff;
s_mem_contents[14'h00e5] = 8'hff;
s_mem_contents[14'h00e6] = 8'hff;
s_mem_contents[14'h00e7] = 8'hff;
s_mem_contents[14'h00e8] = 8'hff;
s_mem_contents[14'h00e9] = 8'hff;
s_mem_contents[14'h00ea] = 8'hff;
s_mem_contents[14'h00eb] = 8'hff;
s_mem_contents[14'h00ec] = 8'hff;
s_mem_contents[14'h00ed] = 8'hff;
s_mem_contents[14'h00ee] = 8'hff;
s_mem_contents[14'h00ef] = 8'hff;
s_mem_contents[14'h00f0] = 8'hff;
s_mem_contents[14'h00f1] = 8'hff;
s_mem_contents[14'h00f2] = 8'hff;
s_mem_contents[14'h00f3] = 8'hff;
s_mem_contents[14'h00f4] = 8'hff;
s_mem_contents[14'h00f5] = 8'hff;
s_mem_contents[14'h00f6] = 8'hff;
s_mem_contents[14'h00f7] = 8'hff;
s_mem_contents[14'h00f8] = 8'hff;
s_mem_contents[14'h00f9] = 8'hff;
s_mem_contents[14'h00fa] = 8'hff;
s_mem_contents[14'h00fb] = 8'hff;
s_mem_contents[14'h00fc] = 8'hff;
s_mem_contents[14'h00fd] = 8'hff;
s_mem_contents[14'h00fe] = 8'hff;
s_mem_contents[14'h00ff] = 8'hff;
s_mem_contents[14'h0100] = 8'hff;
s_mem_contents[14'h0101] = 8'hff;
s_mem_contents[14'h0102] = 8'hff;
s_mem_contents[14'h0103] = 8'hff;
s_mem_contents[14'h0104] = 8'hff;
s_mem_contents[14'h0105] = 8'hff;
s_mem_contents[14'h0106] = 8'hff;
s_mem_contents[14'h0107] = 8'hff;
s_mem_contents[14'h0108] = 8'hff;
s_mem_contents[14'h0109] = 8'hff;
s_mem_contents[14'h010a] = 8'hff;
s_mem_contents[14'h010b] = 8'hff;
s_mem_contents[14'h010c] = 8'hff;
s_mem_contents[14'h010d] = 8'hff;
s_mem_contents[14'h010e] = 8'hff;
s_mem_contents[14'h010f] = 8'hff;
s_mem_contents[14'h0110] = 8'hff;
s_mem_contents[14'h0111] = 8'hff;
s_mem_contents[14'h0112] = 8'hff;
s_mem_contents[14'h0113] = 8'hff;
s_mem_contents[14'h0114] = 8'hff;
s_mem_contents[14'h0115] = 8'hff;
s_mem_contents[14'h0116] = 8'hff;
s_mem_contents[14'h0117] = 8'hff;
s_mem_contents[14'h0118] = 8'hff;
s_mem_contents[14'h0119] = 8'hff;
s_mem_contents[14'h011a] = 8'hff;
s_mem_contents[14'h011b] = 8'hff;
s_mem_contents[14'h011c] = 8'hff;
s_mem_contents[14'h011d] = 8'hff;
s_mem_contents[14'h011e] = 8'hff;
s_mem_contents[14'h011f] = 8'hff;
s_mem_contents[14'h0120] = 8'hff;
s_mem_contents[14'h0121] = 8'hff;
s_mem_contents[14'h0122] = 8'hff;
s_mem_contents[14'h0123] = 8'hff;
s_mem_contents[14'h0124] = 8'hff;
s_mem_contents[14'h0125] = 8'hff;
s_mem_contents[14'h0126] = 8'hff;
s_mem_contents[14'h0127] = 8'hff;
s_mem_contents[14'h0128] = 8'hff;
s_mem_contents[14'h0129] = 8'hff;
s_mem_contents[14'h012a] = 8'hff;
s_mem_contents[14'h012b] = 8'hff;
s_mem_contents[14'h012c] = 8'hff;
s_mem_contents[14'h012d] = 8'hff;
s_mem_contents[14'h012e] = 8'hff;
s_mem_contents[14'h012f] = 8'hff;
s_mem_contents[14'h0130] = 8'hff;
s_mem_contents[14'h0131] = 8'hff;
s_mem_contents[14'h0132] = 8'hff;
s_mem_contents[14'h0133] = 8'hff;
s_mem_contents[14'h0134] = 8'hff;
s_mem_contents[14'h0135] = 8'hff;
s_mem_contents[14'h0136] = 8'hff;
s_mem_contents[14'h0137] = 8'hff;
s_mem_contents[14'h0138] = 8'hff;
s_mem_contents[14'h0139] = 8'hff;
s_mem_contents[14'h013a] = 8'hff;
s_mem_contents[14'h013b] = 8'hff;
s_mem_contents[14'h013c] = 8'hff;
s_mem_contents[14'h013d] = 8'hff;
s_mem_contents[14'h013e] = 8'hff;
s_mem_contents[14'h013f] = 8'hff;
s_mem_contents[14'h0140] = 8'hff;
s_mem_contents[14'h0141] = 8'hff;
s_mem_contents[14'h0142] = 8'hff;
s_mem_contents[14'h0143] = 8'hff;
s_mem_contents[14'h0144] = 8'hff;
s_mem_contents[14'h0145] = 8'hff;
s_mem_contents[14'h0146] = 8'hff;
s_mem_contents[14'h0147] = 8'hff;
s_mem_contents[14'h0148] = 8'hff;
s_mem_contents[14'h0149] = 8'hff;
s_mem_contents[14'h014a] = 8'hff;
s_mem_contents[14'h014b] = 8'hff;
s_mem_contents[14'h014c] = 8'hff;
s_mem_contents[14'h014d] = 8'hff;
s_mem_contents[14'h014e] = 8'hff;
s_mem_contents[14'h014f] = 8'hff;
s_mem_contents[14'h0150] = 8'hff;
s_mem_contents[14'h0151] = 8'hff;
s_mem_contents[14'h0152] = 8'hff;
s_mem_contents[14'h0153] = 8'hff;
s_mem_contents[14'h0154] = 8'hff;
s_mem_contents[14'h0155] = 8'hff;
s_mem_contents[14'h0156] = 8'hff;
s_mem_contents[14'h0157] = 8'hff;
s_mem_contents[14'h0158] = 8'hff;
s_mem_contents[14'h0159] = 8'hff;
s_mem_contents[14'h015a] = 8'hff;
s_mem_contents[14'h015b] = 8'hff;
s_mem_contents[14'h015c] = 8'hff;
s_mem_contents[14'h015d] = 8'hff;
s_mem_contents[14'h015e] = 8'hff;
s_mem_contents[14'h015f] = 8'hff;
s_mem_contents[14'h0160] = 8'hff;
s_mem_contents[14'h0161] = 8'hff;
s_mem_contents[14'h0162] = 8'hff;
s_mem_contents[14'h0163] = 8'hff;
s_mem_contents[14'h0164] = 8'hff;
s_mem_contents[14'h0165] = 8'hff;
s_mem_contents[14'h0166] = 8'hff;
s_mem_contents[14'h0167] = 8'hff;
s_mem_contents[14'h0168] = 8'hff;
s_mem_contents[14'h0169] = 8'hff;
s_mem_contents[14'h016a] = 8'hff;
s_mem_contents[14'h016b] = 8'hff;
s_mem_contents[14'h016c] = 8'hff;
s_mem_contents[14'h016d] = 8'hff;
s_mem_contents[14'h016e] = 8'hff;
s_mem_contents[14'h016f] = 8'hff;
s_mem_contents[14'h0170] = 8'hff;
s_mem_contents[14'h0171] = 8'hff;
s_mem_contents[14'h0172] = 8'hff;
s_mem_contents[14'h0173] = 8'hff;
s_mem_contents[14'h0174] = 8'hff;
s_mem_contents[14'h0175] = 8'hff;
s_mem_contents[14'h0176] = 8'hff;
s_mem_contents[14'h0177] = 8'hff;
s_mem_contents[14'h0178] = 8'hff;
s_mem_contents[14'h0179] = 8'hff;
s_mem_contents[14'h017a] = 8'hff;
s_mem_contents[14'h017b] = 8'hff;
s_mem_contents[14'h017c] = 8'hff;
s_mem_contents[14'h017d] = 8'hff;
s_mem_contents[14'h017e] = 8'hff;
s_mem_contents[14'h017f] = 8'hff;
s_mem_contents[14'h0180] = 8'hff;
s_mem_contents[14'h0181] = 8'hff;
s_mem_contents[14'h0182] = 8'hff;
s_mem_contents[14'h0183] = 8'hff;
s_mem_contents[14'h0184] = 8'hff;
s_mem_contents[14'h0185] = 8'hff;
s_mem_contents[14'h0186] = 8'hff;
s_mem_contents[14'h0187] = 8'hff;
s_mem_contents[14'h0188] = 8'hff;
s_mem_contents[14'h0189] = 8'hff;
s_mem_contents[14'h018a] = 8'hff;
s_mem_contents[14'h018b] = 8'hff;
s_mem_contents[14'h018c] = 8'hff;
s_mem_contents[14'h018d] = 8'hff;
s_mem_contents[14'h018e] = 8'hff;
s_mem_contents[14'h018f] = 8'hff;
s_mem_contents[14'h0190] = 8'hff;
s_mem_contents[14'h0191] = 8'hff;
s_mem_contents[14'h0192] = 8'hff;
s_mem_contents[14'h0193] = 8'hff;
s_mem_contents[14'h0194] = 8'hff;
s_mem_contents[14'h0195] = 8'hff;
s_mem_contents[14'h0196] = 8'hff;
s_mem_contents[14'h0197] = 8'hff;
s_mem_contents[14'h0198] = 8'hff;
s_mem_contents[14'h0199] = 8'hff;
s_mem_contents[14'h019a] = 8'hff;
s_mem_contents[14'h019b] = 8'hff;
s_mem_contents[14'h019c] = 8'hff;
s_mem_contents[14'h019d] = 8'hff;
s_mem_contents[14'h019e] = 8'hff;
s_mem_contents[14'h019f] = 8'hff;
s_mem_contents[14'h01a0] = 8'hff;
s_mem_contents[14'h01a1] = 8'hff;
s_mem_contents[14'h01a2] = 8'hff;
s_mem_contents[14'h01a3] = 8'hff;
s_mem_contents[14'h01a4] = 8'hff;
s_mem_contents[14'h01a5] = 8'hff;
s_mem_contents[14'h01a6] = 8'hff;
s_mem_contents[14'h01a7] = 8'hff;
s_mem_contents[14'h01a8] = 8'hff;
s_mem_contents[14'h01a9] = 8'hff;
s_mem_contents[14'h01aa] = 8'hff;
s_mem_contents[14'h01ab] = 8'hff;
s_mem_contents[14'h01ac] = 8'hff;
s_mem_contents[14'h01ad] = 8'hff;
s_mem_contents[14'h01ae] = 8'hff;
s_mem_contents[14'h01af] = 8'hff;
s_mem_contents[14'h01b0] = 8'hff;
s_mem_contents[14'h01b1] = 8'hff;
s_mem_contents[14'h01b2] = 8'hff;
s_mem_contents[14'h01b3] = 8'hff;
s_mem_contents[14'h01b4] = 8'hff;
s_mem_contents[14'h01b5] = 8'hff;
s_mem_contents[14'h01b6] = 8'hff;
s_mem_contents[14'h01b7] = 8'hff;
s_mem_contents[14'h01b8] = 8'hff;
s_mem_contents[14'h01b9] = 8'hff;
s_mem_contents[14'h01ba] = 8'hff;
s_mem_contents[14'h01bb] = 8'hff;
s_mem_contents[14'h01bc] = 8'hff;
s_mem_contents[14'h01bd] = 8'hff;
s_mem_contents[14'h01be] = 8'hff;
s_mem_contents[14'h01bf] = 8'hff;
s_mem_contents[14'h01c0] = 8'hff;
s_mem_contents[14'h01c1] = 8'hff;
s_mem_contents[14'h01c2] = 8'hff;
s_mem_contents[14'h01c3] = 8'hff;
s_mem_contents[14'h01c4] = 8'hff;
s_mem_contents[14'h01c5] = 8'hff;
s_mem_contents[14'h01c6] = 8'hff;
s_mem_contents[14'h01c7] = 8'hff;
s_mem_contents[14'h01c8] = 8'hff;
s_mem_contents[14'h01c9] = 8'hff;
s_mem_contents[14'h01ca] = 8'hff;
s_mem_contents[14'h01cb] = 8'hff;
s_mem_contents[14'h01cc] = 8'hff;
s_mem_contents[14'h01cd] = 8'hff;
s_mem_contents[14'h01ce] = 8'hff;
s_mem_contents[14'h01cf] = 8'hff;
s_mem_contents[14'h01d0] = 8'hff;
s_mem_contents[14'h01d1] = 8'hff;
s_mem_contents[14'h01d2] = 8'hff;
s_mem_contents[14'h01d3] = 8'hff;
s_mem_contents[14'h01d4] = 8'hff;
s_mem_contents[14'h01d5] = 8'hff;
s_mem_contents[14'h01d6] = 8'hff;
s_mem_contents[14'h01d7] = 8'hff;
s_mem_contents[14'h01d8] = 8'hff;
s_mem_contents[14'h01d9] = 8'hff;
s_mem_contents[14'h01da] = 8'hff;
s_mem_contents[14'h01db] = 8'hff;
s_mem_contents[14'h01dc] = 8'hff;
s_mem_contents[14'h01dd] = 8'hff;
s_mem_contents[14'h01de] = 8'hff;
s_mem_contents[14'h01df] = 8'hff;
s_mem_contents[14'h01e0] = 8'hff;
s_mem_contents[14'h01e1] = 8'hff;
s_mem_contents[14'h01e2] = 8'hff;
s_mem_contents[14'h01e3] = 8'hff;
s_mem_contents[14'h01e4] = 8'hff;
s_mem_contents[14'h01e5] = 8'hff;
s_mem_contents[14'h01e6] = 8'hff;
s_mem_contents[14'h01e7] = 8'hff;
s_mem_contents[14'h01e8] = 8'hff;
s_mem_contents[14'h01e9] = 8'hff;
s_mem_contents[14'h01ea] = 8'hff;
s_mem_contents[14'h01eb] = 8'hff;
s_mem_contents[14'h01ec] = 8'hff;
s_mem_contents[14'h01ed] = 8'hff;
s_mem_contents[14'h01ee] = 8'hff;
s_mem_contents[14'h01ef] = 8'hff;
s_mem_contents[14'h01f0] = 8'hff;
s_mem_contents[14'h01f1] = 8'hff;
s_mem_contents[14'h01f2] = 8'hff;
s_mem_contents[14'h01f3] = 8'hff;
s_mem_contents[14'h01f4] = 8'hff;
s_mem_contents[14'h01f5] = 8'hff;
s_mem_contents[14'h01f6] = 8'hff;
s_mem_contents[14'h01f7] = 8'hff;
s_mem_contents[14'h01f8] = 8'hff;
s_mem_contents[14'h01f9] = 8'hff;
s_mem_contents[14'h01fa] = 8'hff;
s_mem_contents[14'h01fb] = 8'hff;
s_mem_contents[14'h01fc] = 8'hff;
s_mem_contents[14'h01fd] = 8'hff;
s_mem_contents[14'h01fe] = 8'hff;
s_mem_contents[14'h01ff] = 8'hff;
s_mem_contents[14'h0200] = 8'h00;
s_mem_contents[14'h0201] = 8'h00;
s_mem_contents[14'h0202] = 8'h00;
s_mem_contents[14'h0203] = 8'h00;
s_mem_contents[14'h0204] = 8'h00;
s_mem_contents[14'h0205] = 8'h00;
s_mem_contents[14'h0206] = 8'h00;
s_mem_contents[14'h0207] = 8'h00;
s_mem_contents[14'h0208] = 8'h29;
s_mem_contents[14'h0209] = 8'h00;
s_mem_contents[14'h020a] = 8'h60;
s_mem_contents[14'h020b] = 8'h49;
s_mem_contents[14'h020c] = 8'h00;
s_mem_contents[14'h020d] = 8'h60;
s_mem_contents[14'h020e] = 8'h09;
s_mem_contents[14'h020f] = 8'h00;
s_mem_contents[14'h0210] = 8'h60;
s_mem_contents[14'h0211] = 8'h69;
s_mem_contents[14'h0212] = 8'h00;
s_mem_contents[14'h0213] = 8'h60;
s_mem_contents[14'h0214] = 8'he9;
s_mem_contents[14'h0215] = 8'h00;
s_mem_contents[14'h0216] = 8'h60;
s_mem_contents[14'h0217] = 8'hc3;
s_mem_contents[14'h0218] = 8'h82;
s_mem_contents[14'h0219] = 8'h41;
s_mem_contents[14'h021a] = 8'h00;
s_mem_contents[14'h021b] = 8'h7f;
s_mem_contents[14'h021c] = 8'h80;
s_mem_contents[14'h021d] = 8'h80;
s_mem_contents[14'h021e] = 8'h00;
s_mem_contents[14'h021f] = 8'h02;
s_mem_contents[14'h0220] = 8'h86;
s_mem_contents[14'h0221] = 8'h04;
s_mem_contents[14'h0222] = 8'h82;
s_mem_contents[14'h0223] = 8'h00;
s_mem_contents[14'h0224] = 8'h87;
s_mem_contents[14'h0225] = 8'h05;
s_mem_contents[14'h0226] = 8'h83;
s_mem_contents[14'h0227] = 8'h01;
s_mem_contents[14'h0228] = 8'h61;
s_mem_contents[14'h0229] = 8'h41;
s_mem_contents[14'h022a] = 8'h20;
s_mem_contents[14'h022b] = 8'h00;
s_mem_contents[14'h022c] = 8'he1;
s_mem_contents[14'h022d] = 8'hc1;
s_mem_contents[14'h022e] = 8'ha0;
s_mem_contents[14'h022f] = 8'h80;
s_mem_contents[14'h0230] = 8'h81;
s_mem_contents[14'h0231] = 8'h01;
s_mem_contents[14'h0232] = 8'h80;
s_mem_contents[14'h0233] = 8'h02;
s_mem_contents[14'h0234] = 8'h81;
s_mem_contents[14'h0235] = 8'h01;
s_mem_contents[14'h0236] = 8'h80;
s_mem_contents[14'h0237] = 8'h00;
s_mem_contents[14'h0238] = 8'h01;
s_mem_contents[14'h0239] = 8'h00;
s_mem_contents[14'h023a] = 8'h01;
s_mem_contents[14'h023b] = 8'h02;
s_mem_contents[14'h023c] = 8'h81;
s_mem_contents[14'h023d] = 8'h80;
s_mem_contents[14'h023e] = 8'h81;
s_mem_contents[14'h023f] = 8'h80;
s_mem_contents[14'h0240] = 8'h7f;
s_mem_contents[14'h0241] = 8'h80;
s_mem_contents[14'h0242] = 8'hff;
s_mem_contents[14'h0243] = 8'h00;
s_mem_contents[14'h0244] = 8'h01;
s_mem_contents[14'h0245] = 8'h00;
s_mem_contents[14'h0246] = 8'h80;
s_mem_contents[14'h0247] = 8'h80;
s_mem_contents[14'h0248] = 8'h02;
s_mem_contents[14'h0249] = 8'h00;
s_mem_contents[14'h024a] = 8'h00;
s_mem_contents[14'h024b] = 8'h1f;
s_mem_contents[14'h024c] = 8'h71;
s_mem_contents[14'h024d] = 8'h80;
s_mem_contents[14'h024e] = 8'h0f;
s_mem_contents[14'h024f] = 8'hff;
s_mem_contents[14'h0250] = 8'h7f;
s_mem_contents[14'h0251] = 8'h80;
s_mem_contents[14'h0252] = 8'hff;
s_mem_contents[14'h0253] = 8'h0f;
s_mem_contents[14'h0254] = 8'h8f;
s_mem_contents[14'h0255] = 8'h8f;
s_mem_contents[14'h0256] = 8'h00;
s_mem_contents[14'h0257] = 8'hf1;
s_mem_contents[14'h0258] = 8'h1f;
s_mem_contents[14'h0259] = 8'h00;
s_mem_contents[14'h025a] = 8'hf0;
s_mem_contents[14'h025b] = 8'hff;
s_mem_contents[14'h025c] = 8'hff;
s_mem_contents[14'h025d] = 8'hff;
s_mem_contents[14'h025e] = 8'hff;
s_mem_contents[14'h025f] = 8'hf0;
s_mem_contents[14'h0260] = 8'hf0;
s_mem_contents[14'h0261] = 8'h0f;
s_mem_contents[14'h0262] = 8'h00;
s_mem_contents[14'h0263] = 8'hff;
s_mem_contents[14'h0264] = 8'h7f;
s_mem_contents[14'h0265] = 8'h80;
s_mem_contents[14'h0266] = 8'h02;
s_mem_contents[14'h0267] = 8'h80;
s_mem_contents[14'h0268] = 8'h00;
s_mem_contents[14'h0269] = 8'h80;
s_mem_contents[14'h026a] = 8'hff;
s_mem_contents[14'h026b] = 8'hff;
s_mem_contents[14'h026c] = 8'hff;
s_mem_contents[14'h026d] = 8'hff;
s_mem_contents[14'h026e] = 8'hff;
s_mem_contents[14'h026f] = 8'hff;
s_mem_contents[14'h0270] = 8'hff;
s_mem_contents[14'h0271] = 8'hff;
s_mem_contents[14'h0272] = 8'hff;
s_mem_contents[14'h0273] = 8'hff;
s_mem_contents[14'h0274] = 8'hff;
s_mem_contents[14'h0275] = 8'hff;
s_mem_contents[14'h0276] = 8'hff;
s_mem_contents[14'h0277] = 8'hff;
s_mem_contents[14'h0278] = 8'hff;
s_mem_contents[14'h0279] = 8'hff;
s_mem_contents[14'h027a] = 8'hff;
s_mem_contents[14'h027b] = 8'hff;
s_mem_contents[14'h027c] = 8'hff;
s_mem_contents[14'h027d] = 8'hff;
s_mem_contents[14'h027e] = 8'hff;
s_mem_contents[14'h027f] = 8'hff;
s_mem_contents[14'h0280] = 8'hff;
s_mem_contents[14'h0281] = 8'hff;
s_mem_contents[14'h0282] = 8'hff;
s_mem_contents[14'h0283] = 8'hff;
s_mem_contents[14'h0284] = 8'hff;
s_mem_contents[14'h0285] = 8'hff;
s_mem_contents[14'h0286] = 8'hff;
s_mem_contents[14'h0287] = 8'hff;
s_mem_contents[14'h0288] = 8'hff;
s_mem_contents[14'h0289] = 8'hff;
s_mem_contents[14'h028a] = 8'hff;
s_mem_contents[14'h028b] = 8'hff;
s_mem_contents[14'h028c] = 8'hff;
s_mem_contents[14'h028d] = 8'hff;
s_mem_contents[14'h028e] = 8'hff;
s_mem_contents[14'h028f] = 8'hff;
s_mem_contents[14'h0290] = 8'hff;
s_mem_contents[14'h0291] = 8'hff;
s_mem_contents[14'h0292] = 8'hff;
s_mem_contents[14'h0293] = 8'hff;
s_mem_contents[14'h0294] = 8'hff;
s_mem_contents[14'h0295] = 8'hff;
s_mem_contents[14'h0296] = 8'hff;
s_mem_contents[14'h0297] = 8'hff;
s_mem_contents[14'h0298] = 8'hff;
s_mem_contents[14'h0299] = 8'hff;
s_mem_contents[14'h029a] = 8'hff;
s_mem_contents[14'h029b] = 8'hff;
s_mem_contents[14'h029c] = 8'hff;
s_mem_contents[14'h029d] = 8'hff;
s_mem_contents[14'h029e] = 8'hff;
s_mem_contents[14'h029f] = 8'hff;
s_mem_contents[14'h02a0] = 8'hff;
s_mem_contents[14'h02a1] = 8'hff;
s_mem_contents[14'h02a2] = 8'hff;
s_mem_contents[14'h02a3] = 8'hff;
s_mem_contents[14'h02a4] = 8'hff;
s_mem_contents[14'h02a5] = 8'hff;
s_mem_contents[14'h02a6] = 8'hff;
s_mem_contents[14'h02a7] = 8'hff;
s_mem_contents[14'h02a8] = 8'hff;
s_mem_contents[14'h02a9] = 8'hff;
s_mem_contents[14'h02aa] = 8'hff;
s_mem_contents[14'h02ab] = 8'hff;
s_mem_contents[14'h02ac] = 8'hff;
s_mem_contents[14'h02ad] = 8'hff;
s_mem_contents[14'h02ae] = 8'hff;
s_mem_contents[14'h02af] = 8'hff;
s_mem_contents[14'h02b0] = 8'hff;
s_mem_contents[14'h02b1] = 8'hff;
s_mem_contents[14'h02b2] = 8'hff;
s_mem_contents[14'h02b3] = 8'hff;
s_mem_contents[14'h02b4] = 8'hff;
s_mem_contents[14'h02b5] = 8'hff;
s_mem_contents[14'h02b6] = 8'hff;
s_mem_contents[14'h02b7] = 8'hff;
s_mem_contents[14'h02b8] = 8'hff;
s_mem_contents[14'h02b9] = 8'hff;
s_mem_contents[14'h02ba] = 8'hff;
s_mem_contents[14'h02bb] = 8'hff;
s_mem_contents[14'h02bc] = 8'hff;
s_mem_contents[14'h02bd] = 8'hff;
s_mem_contents[14'h02be] = 8'hff;
s_mem_contents[14'h02bf] = 8'hff;
s_mem_contents[14'h02c0] = 8'hff;
s_mem_contents[14'h02c1] = 8'hff;
s_mem_contents[14'h02c2] = 8'hff;
s_mem_contents[14'h02c3] = 8'hff;
s_mem_contents[14'h02c4] = 8'hff;
s_mem_contents[14'h02c5] = 8'hff;
s_mem_contents[14'h02c6] = 8'hff;
s_mem_contents[14'h02c7] = 8'hff;
s_mem_contents[14'h02c8] = 8'hff;
s_mem_contents[14'h02c9] = 8'hff;
s_mem_contents[14'h02ca] = 8'hff;
s_mem_contents[14'h02cb] = 8'hff;
s_mem_contents[14'h02cc] = 8'hff;
s_mem_contents[14'h02cd] = 8'hff;
s_mem_contents[14'h02ce] = 8'hff;
s_mem_contents[14'h02cf] = 8'hff;
s_mem_contents[14'h02d0] = 8'hff;
s_mem_contents[14'h02d1] = 8'hff;
s_mem_contents[14'h02d2] = 8'hff;
s_mem_contents[14'h02d3] = 8'hff;
s_mem_contents[14'h02d4] = 8'hff;
s_mem_contents[14'h02d5] = 8'hff;
s_mem_contents[14'h02d6] = 8'hff;
s_mem_contents[14'h02d7] = 8'hff;
s_mem_contents[14'h02d8] = 8'hff;
s_mem_contents[14'h02d9] = 8'hff;
s_mem_contents[14'h02da] = 8'hff;
s_mem_contents[14'h02db] = 8'hff;
s_mem_contents[14'h02dc] = 8'hff;
s_mem_contents[14'h02dd] = 8'hff;
s_mem_contents[14'h02de] = 8'hff;
s_mem_contents[14'h02df] = 8'hff;
s_mem_contents[14'h02e0] = 8'hff;
s_mem_contents[14'h02e1] = 8'hff;
s_mem_contents[14'h02e2] = 8'hff;
s_mem_contents[14'h02e3] = 8'hff;
s_mem_contents[14'h02e4] = 8'hff;
s_mem_contents[14'h02e5] = 8'hff;
s_mem_contents[14'h02e6] = 8'hff;
s_mem_contents[14'h02e7] = 8'hff;
s_mem_contents[14'h02e8] = 8'hff;
s_mem_contents[14'h02e9] = 8'hff;
s_mem_contents[14'h02ea] = 8'hff;
s_mem_contents[14'h02eb] = 8'hff;
s_mem_contents[14'h02ec] = 8'hff;
s_mem_contents[14'h02ed] = 8'hff;
s_mem_contents[14'h02ee] = 8'hff;
s_mem_contents[14'h02ef] = 8'hff;
s_mem_contents[14'h02f0] = 8'hff;
s_mem_contents[14'h02f1] = 8'hff;
s_mem_contents[14'h02f2] = 8'hff;
s_mem_contents[14'h02f3] = 8'hff;
s_mem_contents[14'h02f4] = 8'hff;
s_mem_contents[14'h02f5] = 8'hff;
s_mem_contents[14'h02f6] = 8'hff;
s_mem_contents[14'h02f7] = 8'hff;
s_mem_contents[14'h02f8] = 8'hff;
s_mem_contents[14'h02f9] = 8'hff;
s_mem_contents[14'h02fa] = 8'hff;
s_mem_contents[14'h02fb] = 8'hff;
s_mem_contents[14'h02fc] = 8'hff;
s_mem_contents[14'h02fd] = 8'hff;
s_mem_contents[14'h02fe] = 8'hff;
s_mem_contents[14'h02ff] = 8'hff;
s_mem_contents[14'h0300] = 8'hff;
s_mem_contents[14'h0301] = 8'hff;
s_mem_contents[14'h0302] = 8'hff;
s_mem_contents[14'h0303] = 8'hff;
s_mem_contents[14'h0304] = 8'hff;
s_mem_contents[14'h0305] = 8'hff;
s_mem_contents[14'h0306] = 8'hff;
s_mem_contents[14'h0307] = 8'hff;
s_mem_contents[14'h0308] = 8'hff;
s_mem_contents[14'h0309] = 8'hff;
s_mem_contents[14'h030a] = 8'hff;
s_mem_contents[14'h030b] = 8'hff;
s_mem_contents[14'h030c] = 8'hff;
s_mem_contents[14'h030d] = 8'hff;
s_mem_contents[14'h030e] = 8'hff;
s_mem_contents[14'h030f] = 8'hff;
s_mem_contents[14'h0310] = 8'hff;
s_mem_contents[14'h0311] = 8'hff;
s_mem_contents[14'h0312] = 8'hff;
s_mem_contents[14'h0313] = 8'hff;
s_mem_contents[14'h0314] = 8'hff;
s_mem_contents[14'h0315] = 8'hff;
s_mem_contents[14'h0316] = 8'hff;
s_mem_contents[14'h0317] = 8'hff;
s_mem_contents[14'h0318] = 8'hff;
s_mem_contents[14'h0319] = 8'hff;
s_mem_contents[14'h031a] = 8'hff;
s_mem_contents[14'h031b] = 8'hff;
s_mem_contents[14'h031c] = 8'hff;
s_mem_contents[14'h031d] = 8'hff;
s_mem_contents[14'h031e] = 8'hff;
s_mem_contents[14'h031f] = 8'hff;
s_mem_contents[14'h0320] = 8'hff;
s_mem_contents[14'h0321] = 8'hff;
s_mem_contents[14'h0322] = 8'hff;
s_mem_contents[14'h0323] = 8'hff;
s_mem_contents[14'h0324] = 8'hff;
s_mem_contents[14'h0325] = 8'hff;
s_mem_contents[14'h0326] = 8'hff;
s_mem_contents[14'h0327] = 8'hff;
s_mem_contents[14'h0328] = 8'hff;
s_mem_contents[14'h0329] = 8'hff;
s_mem_contents[14'h032a] = 8'hff;
s_mem_contents[14'h032b] = 8'hff;
s_mem_contents[14'h032c] = 8'hff;
s_mem_contents[14'h032d] = 8'hff;
s_mem_contents[14'h032e] = 8'hff;
s_mem_contents[14'h032f] = 8'hff;
s_mem_contents[14'h0330] = 8'hff;
s_mem_contents[14'h0331] = 8'hff;
s_mem_contents[14'h0332] = 8'hff;
s_mem_contents[14'h0333] = 8'hff;
s_mem_contents[14'h0334] = 8'hff;
s_mem_contents[14'h0335] = 8'hff;
s_mem_contents[14'h0336] = 8'hff;
s_mem_contents[14'h0337] = 8'hff;
s_mem_contents[14'h0338] = 8'hff;
s_mem_contents[14'h0339] = 8'hff;
s_mem_contents[14'h033a] = 8'hff;
s_mem_contents[14'h033b] = 8'hff;
s_mem_contents[14'h033c] = 8'hff;
s_mem_contents[14'h033d] = 8'hff;
s_mem_contents[14'h033e] = 8'hff;
s_mem_contents[14'h033f] = 8'hff;
s_mem_contents[14'h0340] = 8'hff;
s_mem_contents[14'h0341] = 8'hff;
s_mem_contents[14'h0342] = 8'hff;
s_mem_contents[14'h0343] = 8'hff;
s_mem_contents[14'h0344] = 8'hff;
s_mem_contents[14'h0345] = 8'hff;
s_mem_contents[14'h0346] = 8'hff;
s_mem_contents[14'h0347] = 8'hff;
s_mem_contents[14'h0348] = 8'hff;
s_mem_contents[14'h0349] = 8'hff;
s_mem_contents[14'h034a] = 8'hff;
s_mem_contents[14'h034b] = 8'hff;
s_mem_contents[14'h034c] = 8'hff;
s_mem_contents[14'h034d] = 8'hff;
s_mem_contents[14'h034e] = 8'hff;
s_mem_contents[14'h034f] = 8'hff;
s_mem_contents[14'h0350] = 8'hff;
s_mem_contents[14'h0351] = 8'hff;
s_mem_contents[14'h0352] = 8'hff;
s_mem_contents[14'h0353] = 8'hff;
s_mem_contents[14'h0354] = 8'hff;
s_mem_contents[14'h0355] = 8'hff;
s_mem_contents[14'h0356] = 8'hff;
s_mem_contents[14'h0357] = 8'hff;
s_mem_contents[14'h0358] = 8'hff;
s_mem_contents[14'h0359] = 8'hff;
s_mem_contents[14'h035a] = 8'hff;
s_mem_contents[14'h035b] = 8'hff;
s_mem_contents[14'h035c] = 8'hff;
s_mem_contents[14'h035d] = 8'hff;
s_mem_contents[14'h035e] = 8'hff;
s_mem_contents[14'h035f] = 8'hff;
s_mem_contents[14'h0360] = 8'hff;
s_mem_contents[14'h0361] = 8'hff;
s_mem_contents[14'h0362] = 8'hff;
s_mem_contents[14'h0363] = 8'hff;
s_mem_contents[14'h0364] = 8'hff;
s_mem_contents[14'h0365] = 8'hff;
s_mem_contents[14'h0366] = 8'hff;
s_mem_contents[14'h0367] = 8'hff;
s_mem_contents[14'h0368] = 8'hff;
s_mem_contents[14'h0369] = 8'hff;
s_mem_contents[14'h036a] = 8'hff;
s_mem_contents[14'h036b] = 8'hff;
s_mem_contents[14'h036c] = 8'hff;
s_mem_contents[14'h036d] = 8'hff;
s_mem_contents[14'h036e] = 8'hff;
s_mem_contents[14'h036f] = 8'hff;
s_mem_contents[14'h0370] = 8'hff;
s_mem_contents[14'h0371] = 8'hff;
s_mem_contents[14'h0372] = 8'hff;
s_mem_contents[14'h0373] = 8'hff;
s_mem_contents[14'h0374] = 8'hff;
s_mem_contents[14'h0375] = 8'hff;
s_mem_contents[14'h0376] = 8'hff;
s_mem_contents[14'h0377] = 8'hff;
s_mem_contents[14'h0378] = 8'hff;
s_mem_contents[14'h0379] = 8'hff;
s_mem_contents[14'h037a] = 8'hff;
s_mem_contents[14'h037b] = 8'hff;
s_mem_contents[14'h037c] = 8'hff;
s_mem_contents[14'h037d] = 8'hff;
s_mem_contents[14'h037e] = 8'hff;
s_mem_contents[14'h037f] = 8'hff;
s_mem_contents[14'h0380] = 8'hff;
s_mem_contents[14'h0381] = 8'hff;
s_mem_contents[14'h0382] = 8'hff;
s_mem_contents[14'h0383] = 8'hff;
s_mem_contents[14'h0384] = 8'hff;
s_mem_contents[14'h0385] = 8'hff;
s_mem_contents[14'h0386] = 8'hff;
s_mem_contents[14'h0387] = 8'hff;
s_mem_contents[14'h0388] = 8'hff;
s_mem_contents[14'h0389] = 8'hff;
s_mem_contents[14'h038a] = 8'hff;
s_mem_contents[14'h038b] = 8'hff;
s_mem_contents[14'h038c] = 8'hff;
s_mem_contents[14'h038d] = 8'hff;
s_mem_contents[14'h038e] = 8'hff;
s_mem_contents[14'h038f] = 8'hff;
s_mem_contents[14'h0390] = 8'hff;
s_mem_contents[14'h0391] = 8'hff;
s_mem_contents[14'h0392] = 8'hff;
s_mem_contents[14'h0393] = 8'hff;
s_mem_contents[14'h0394] = 8'hff;
s_mem_contents[14'h0395] = 8'hff;
s_mem_contents[14'h0396] = 8'hff;
s_mem_contents[14'h0397] = 8'hff;
s_mem_contents[14'h0398] = 8'hff;
s_mem_contents[14'h0399] = 8'hff;
s_mem_contents[14'h039a] = 8'hff;
s_mem_contents[14'h039b] = 8'hff;
s_mem_contents[14'h039c] = 8'hff;
s_mem_contents[14'h039d] = 8'hff;
s_mem_contents[14'h039e] = 8'hff;
s_mem_contents[14'h039f] = 8'hff;
s_mem_contents[14'h03a0] = 8'hff;
s_mem_contents[14'h03a1] = 8'hff;
s_mem_contents[14'h03a2] = 8'hff;
s_mem_contents[14'h03a3] = 8'hff;
s_mem_contents[14'h03a4] = 8'hff;
s_mem_contents[14'h03a5] = 8'hff;
s_mem_contents[14'h03a6] = 8'hff;
s_mem_contents[14'h03a7] = 8'hff;
s_mem_contents[14'h03a8] = 8'hff;
s_mem_contents[14'h03a9] = 8'hff;
s_mem_contents[14'h03aa] = 8'hff;
s_mem_contents[14'h03ab] = 8'hff;
s_mem_contents[14'h03ac] = 8'hff;
s_mem_contents[14'h03ad] = 8'hff;
s_mem_contents[14'h03ae] = 8'hff;
s_mem_contents[14'h03af] = 8'hff;
s_mem_contents[14'h03b0] = 8'hff;
s_mem_contents[14'h03b1] = 8'hff;
s_mem_contents[14'h03b2] = 8'hff;
s_mem_contents[14'h03b3] = 8'hff;
s_mem_contents[14'h03b4] = 8'hff;
s_mem_contents[14'h03b5] = 8'hff;
s_mem_contents[14'h03b6] = 8'hff;
s_mem_contents[14'h03b7] = 8'hff;
s_mem_contents[14'h03b8] = 8'hff;
s_mem_contents[14'h03b9] = 8'hff;
s_mem_contents[14'h03ba] = 8'hff;
s_mem_contents[14'h03bb] = 8'hff;
s_mem_contents[14'h03bc] = 8'hff;
s_mem_contents[14'h03bd] = 8'hff;
s_mem_contents[14'h03be] = 8'hff;
s_mem_contents[14'h03bf] = 8'hff;
s_mem_contents[14'h03c0] = 8'hff;
s_mem_contents[14'h03c1] = 8'hff;
s_mem_contents[14'h03c2] = 8'hff;
s_mem_contents[14'h03c3] = 8'hff;
s_mem_contents[14'h03c4] = 8'hff;
s_mem_contents[14'h03c5] = 8'hff;
s_mem_contents[14'h03c6] = 8'hff;
s_mem_contents[14'h03c7] = 8'hff;
s_mem_contents[14'h03c8] = 8'hff;
s_mem_contents[14'h03c9] = 8'hff;
s_mem_contents[14'h03ca] = 8'hff;
s_mem_contents[14'h03cb] = 8'hff;
s_mem_contents[14'h03cc] = 8'hff;
s_mem_contents[14'h03cd] = 8'hff;
s_mem_contents[14'h03ce] = 8'hff;
s_mem_contents[14'h03cf] = 8'hff;
s_mem_contents[14'h03d0] = 8'hff;
s_mem_contents[14'h03d1] = 8'hff;
s_mem_contents[14'h03d2] = 8'hff;
s_mem_contents[14'h03d3] = 8'hff;
s_mem_contents[14'h03d4] = 8'hff;
s_mem_contents[14'h03d5] = 8'hff;
s_mem_contents[14'h03d6] = 8'hff;
s_mem_contents[14'h03d7] = 8'hff;
s_mem_contents[14'h03d8] = 8'hff;
s_mem_contents[14'h03d9] = 8'hff;
s_mem_contents[14'h03da] = 8'hff;
s_mem_contents[14'h03db] = 8'hff;
s_mem_contents[14'h03dc] = 8'hff;
s_mem_contents[14'h03dd] = 8'hff;
s_mem_contents[14'h03de] = 8'hff;
s_mem_contents[14'h03df] = 8'hff;
s_mem_contents[14'h03e0] = 8'hff;
s_mem_contents[14'h03e1] = 8'hff;
s_mem_contents[14'h03e2] = 8'hff;
s_mem_contents[14'h03e3] = 8'hff;
s_mem_contents[14'h03e4] = 8'hff;
s_mem_contents[14'h03e5] = 8'hff;
s_mem_contents[14'h03e6] = 8'hff;
s_mem_contents[14'h03e7] = 8'hff;
s_mem_contents[14'h03e8] = 8'hff;
s_mem_contents[14'h03e9] = 8'hff;
s_mem_contents[14'h03ea] = 8'hff;
s_mem_contents[14'h03eb] = 8'hff;
s_mem_contents[14'h03ec] = 8'hff;
s_mem_contents[14'h03ed] = 8'hff;
s_mem_contents[14'h03ee] = 8'hff;
s_mem_contents[14'h03ef] = 8'hff;
s_mem_contents[14'h03f0] = 8'hff;
s_mem_contents[14'h03f1] = 8'hff;
s_mem_contents[14'h03f2] = 8'hff;
s_mem_contents[14'h03f3] = 8'hff;
s_mem_contents[14'h03f4] = 8'hff;
s_mem_contents[14'h03f5] = 8'hff;
s_mem_contents[14'h03f6] = 8'hff;
s_mem_contents[14'h03f7] = 8'hff;
s_mem_contents[14'h03f8] = 8'hff;
s_mem_contents[14'h03f9] = 8'hff;
s_mem_contents[14'h03fa] = 8'hff;
s_mem_contents[14'h03fb] = 8'hff;
s_mem_contents[14'h03fc] = 8'hff;
s_mem_contents[14'h03fd] = 8'hff;
s_mem_contents[14'h03fe] = 8'hff;
s_mem_contents[14'h03ff] = 8'hff;
s_mem_contents[14'h0400] = 8'hd8;
s_mem_contents[14'h0401] = 8'ha2;
s_mem_contents[14'h0402] = 8'hff;
s_mem_contents[14'h0403] = 8'h9a;
s_mem_contents[14'h0404] = 8'ha9;
s_mem_contents[14'h0405] = 8'h00;
s_mem_contents[14'h0406] = 8'h8d;
s_mem_contents[14'h0407] = 8'h00;
s_mem_contents[14'h0408] = 8'h02;
s_mem_contents[14'h0409] = 8'ha2;
s_mem_contents[14'h040a] = 8'h05;
s_mem_contents[14'h040b] = 8'h4c;
s_mem_contents[14'h040c] = 8'h33;
s_mem_contents[14'h040d] = 8'h04;
s_mem_contents[14'h040e] = 8'ha0;
s_mem_contents[14'h040f] = 8'h05;
s_mem_contents[14'h0410] = 8'hd0;
s_mem_contents[14'h0411] = 8'h08;
s_mem_contents[14'h0412] = 8'h4c;
s_mem_contents[14'h0413] = 8'h12;
s_mem_contents[14'h0414] = 8'h04;
s_mem_contents[14'h0415] = 8'h88;
s_mem_contents[14'h0416] = 8'h88;
s_mem_contents[14'h0417] = 8'h88;
s_mem_contents[14'h0418] = 8'h88;
s_mem_contents[14'h0419] = 8'h88;
s_mem_contents[14'h041a] = 8'h88;
s_mem_contents[14'h041b] = 8'h88;
s_mem_contents[14'h041c] = 8'h88;
s_mem_contents[14'h041d] = 8'h88;
s_mem_contents[14'h041e] = 8'h88;
s_mem_contents[14'h041f] = 8'hf0;
s_mem_contents[14'h0420] = 8'h17;
s_mem_contents[14'h0421] = 8'h4c;
s_mem_contents[14'h0422] = 8'h21;
s_mem_contents[14'h0423] = 8'h04;
s_mem_contents[14'h0424] = 8'hca;
s_mem_contents[14'h0425] = 8'hca;
s_mem_contents[14'h0426] = 8'hca;
s_mem_contents[14'h0427] = 8'hca;
s_mem_contents[14'h0428] = 8'hca;
s_mem_contents[14'h0429] = 8'hca;
s_mem_contents[14'h042a] = 8'hca;
s_mem_contents[14'h042b] = 8'hca;
s_mem_contents[14'h042c] = 8'hca;
s_mem_contents[14'h042d] = 8'hca;
s_mem_contents[14'h042e] = 8'hf0;
s_mem_contents[14'h042f] = 8'hde;
s_mem_contents[14'h0430] = 8'h4c;
s_mem_contents[14'h0431] = 8'h30;
s_mem_contents[14'h0432] = 8'h04;
s_mem_contents[14'h0433] = 8'hd0;
s_mem_contents[14'h0434] = 8'hf4;
s_mem_contents[14'h0435] = 8'h4c;
s_mem_contents[14'h0436] = 8'h35;
s_mem_contents[14'h0437] = 8'h04;
s_mem_contents[14'h0438] = 8'had;
s_mem_contents[14'h0439] = 8'h00;
s_mem_contents[14'h043a] = 8'h02;
s_mem_contents[14'h043b] = 8'hc9;
s_mem_contents[14'h043c] = 8'h00;
s_mem_contents[14'h043d] = 8'hd0;
s_mem_contents[14'h043e] = 8'hfe;
s_mem_contents[14'h043f] = 8'ha9;
s_mem_contents[14'h0440] = 8'h01;
s_mem_contents[14'h0441] = 8'h8d;
s_mem_contents[14'h0442] = 8'h00;
s_mem_contents[14'h0443] = 8'h02;
s_mem_contents[14'h0444] = 8'ha0;
s_mem_contents[14'h0445] = 8'hfe;
s_mem_contents[14'h0446] = 8'h88;
s_mem_contents[14'h0447] = 8'h98;
s_mem_contents[14'h0448] = 8'haa;
s_mem_contents[14'h0449] = 8'h10;
s_mem_contents[14'h044a] = 8'h08;
s_mem_contents[14'h044b] = 8'h18;
s_mem_contents[14'h044c] = 8'h69;
s_mem_contents[14'h044d] = 8'h02;
s_mem_contents[14'h044e] = 8'hea;
s_mem_contents[14'h044f] = 8'hea;
s_mem_contents[14'h0450] = 8'hea;
s_mem_contents[14'h0451] = 8'hea;
s_mem_contents[14'h0452] = 8'hea;
s_mem_contents[14'h0453] = 8'hea;
s_mem_contents[14'h0454] = 8'hea;
s_mem_contents[14'h0455] = 8'hea;
s_mem_contents[14'h0456] = 8'hea;
s_mem_contents[14'h0457] = 8'hea;
s_mem_contents[14'h0458] = 8'h49;
s_mem_contents[14'h0459] = 8'h7f;
s_mem_contents[14'h045a] = 8'h8d;
s_mem_contents[14'h045b] = 8'he6;
s_mem_contents[14'h045c] = 8'h04;
s_mem_contents[14'h045d] = 8'ha9;
s_mem_contents[14'h045e] = 8'h00;
s_mem_contents[14'h045f] = 8'h4c;
s_mem_contents[14'h0460] = 8'he5;
s_mem_contents[14'h0461] = 8'h04;
s_mem_contents[14'h0462] = 8'hca;
s_mem_contents[14'h0463] = 8'hca;
s_mem_contents[14'h0464] = 8'hca;
s_mem_contents[14'h0465] = 8'hca;
s_mem_contents[14'h0466] = 8'hca;
s_mem_contents[14'h0467] = 8'hca;
s_mem_contents[14'h0468] = 8'hca;
s_mem_contents[14'h0469] = 8'hca;
s_mem_contents[14'h046a] = 8'hca;
s_mem_contents[14'h046b] = 8'hca;
s_mem_contents[14'h046c] = 8'hca;
s_mem_contents[14'h046d] = 8'hca;
s_mem_contents[14'h046e] = 8'hca;
s_mem_contents[14'h046f] = 8'hca;
s_mem_contents[14'h0470] = 8'hca;
s_mem_contents[14'h0471] = 8'hca;
s_mem_contents[14'h0472] = 8'hca;
s_mem_contents[14'h0473] = 8'hca;
s_mem_contents[14'h0474] = 8'hca;
s_mem_contents[14'h0475] = 8'hca;
s_mem_contents[14'h0476] = 8'hca;
s_mem_contents[14'h0477] = 8'hca;
s_mem_contents[14'h0478] = 8'hca;
s_mem_contents[14'h0479] = 8'hca;
s_mem_contents[14'h047a] = 8'hca;
s_mem_contents[14'h047b] = 8'hca;
s_mem_contents[14'h047c] = 8'hca;
s_mem_contents[14'h047d] = 8'hca;
s_mem_contents[14'h047e] = 8'hca;
s_mem_contents[14'h047f] = 8'hca;
s_mem_contents[14'h0480] = 8'hca;
s_mem_contents[14'h0481] = 8'hca;
s_mem_contents[14'h0482] = 8'hca;
s_mem_contents[14'h0483] = 8'hca;
s_mem_contents[14'h0484] = 8'hca;
s_mem_contents[14'h0485] = 8'hca;
s_mem_contents[14'h0486] = 8'hca;
s_mem_contents[14'h0487] = 8'hca;
s_mem_contents[14'h0488] = 8'hca;
s_mem_contents[14'h0489] = 8'hca;
s_mem_contents[14'h048a] = 8'hca;
s_mem_contents[14'h048b] = 8'hca;
s_mem_contents[14'h048c] = 8'hca;
s_mem_contents[14'h048d] = 8'hca;
s_mem_contents[14'h048e] = 8'hca;
s_mem_contents[14'h048f] = 8'hca;
s_mem_contents[14'h0490] = 8'hca;
s_mem_contents[14'h0491] = 8'hca;
s_mem_contents[14'h0492] = 8'hca;
s_mem_contents[14'h0493] = 8'hca;
s_mem_contents[14'h0494] = 8'hca;
s_mem_contents[14'h0495] = 8'hca;
s_mem_contents[14'h0496] = 8'hca;
s_mem_contents[14'h0497] = 8'hca;
s_mem_contents[14'h0498] = 8'hca;
s_mem_contents[14'h0499] = 8'hca;
s_mem_contents[14'h049a] = 8'hca;
s_mem_contents[14'h049b] = 8'hca;
s_mem_contents[14'h049c] = 8'hca;
s_mem_contents[14'h049d] = 8'hca;
s_mem_contents[14'h049e] = 8'hca;
s_mem_contents[14'h049f] = 8'hca;
s_mem_contents[14'h04a0] = 8'hca;
s_mem_contents[14'h04a1] = 8'hca;
s_mem_contents[14'h04a2] = 8'hca;
s_mem_contents[14'h04a3] = 8'hca;
s_mem_contents[14'h04a4] = 8'hca;
s_mem_contents[14'h04a5] = 8'hca;
s_mem_contents[14'h04a6] = 8'hca;
s_mem_contents[14'h04a7] = 8'hca;
s_mem_contents[14'h04a8] = 8'hca;
s_mem_contents[14'h04a9] = 8'hca;
s_mem_contents[14'h04aa] = 8'hca;
s_mem_contents[14'h04ab] = 8'hca;
s_mem_contents[14'h04ac] = 8'hca;
s_mem_contents[14'h04ad] = 8'hca;
s_mem_contents[14'h04ae] = 8'hca;
s_mem_contents[14'h04af] = 8'hca;
s_mem_contents[14'h04b0] = 8'hca;
s_mem_contents[14'h04b1] = 8'hca;
s_mem_contents[14'h04b2] = 8'hca;
s_mem_contents[14'h04b3] = 8'hca;
s_mem_contents[14'h04b4] = 8'hca;
s_mem_contents[14'h04b5] = 8'hca;
s_mem_contents[14'h04b6] = 8'hca;
s_mem_contents[14'h04b7] = 8'hca;
s_mem_contents[14'h04b8] = 8'hca;
s_mem_contents[14'h04b9] = 8'hca;
s_mem_contents[14'h04ba] = 8'hca;
s_mem_contents[14'h04bb] = 8'hca;
s_mem_contents[14'h04bc] = 8'hca;
s_mem_contents[14'h04bd] = 8'hca;
s_mem_contents[14'h04be] = 8'hca;
s_mem_contents[14'h04bf] = 8'hca;
s_mem_contents[14'h04c0] = 8'hca;
s_mem_contents[14'h04c1] = 8'hca;
s_mem_contents[14'h04c2] = 8'hca;
s_mem_contents[14'h04c3] = 8'hca;
s_mem_contents[14'h04c4] = 8'hca;
s_mem_contents[14'h04c5] = 8'hca;
s_mem_contents[14'h04c6] = 8'hca;
s_mem_contents[14'h04c7] = 8'hca;
s_mem_contents[14'h04c8] = 8'hca;
s_mem_contents[14'h04c9] = 8'hca;
s_mem_contents[14'h04ca] = 8'hca;
s_mem_contents[14'h04cb] = 8'hca;
s_mem_contents[14'h04cc] = 8'hca;
s_mem_contents[14'h04cd] = 8'hca;
s_mem_contents[14'h04ce] = 8'hca;
s_mem_contents[14'h04cf] = 8'hca;
s_mem_contents[14'h04d0] = 8'hca;
s_mem_contents[14'h04d1] = 8'hca;
s_mem_contents[14'h04d2] = 8'hca;
s_mem_contents[14'h04d3] = 8'hca;
s_mem_contents[14'h04d4] = 8'hca;
s_mem_contents[14'h04d5] = 8'hca;
s_mem_contents[14'h04d6] = 8'hca;
s_mem_contents[14'h04d7] = 8'hca;
s_mem_contents[14'h04d8] = 8'hca;
s_mem_contents[14'h04d9] = 8'hca;
s_mem_contents[14'h04da] = 8'hca;
s_mem_contents[14'h04db] = 8'hca;
s_mem_contents[14'h04dc] = 8'hca;
s_mem_contents[14'h04dd] = 8'hca;
s_mem_contents[14'h04de] = 8'hca;
s_mem_contents[14'h04df] = 8'hca;
s_mem_contents[14'h04e0] = 8'hca;
s_mem_contents[14'h04e1] = 8'hca;
s_mem_contents[14'h04e2] = 8'hca;
s_mem_contents[14'h04e3] = 8'hca;
s_mem_contents[14'h04e4] = 8'hca;
s_mem_contents[14'h04e5] = 8'hf0;
s_mem_contents[14'h04e6] = 8'h3e;
s_mem_contents[14'h04e7] = 8'hca;
s_mem_contents[14'h04e8] = 8'hca;
s_mem_contents[14'h04e9] = 8'hca;
s_mem_contents[14'h04ea] = 8'hca;
s_mem_contents[14'h04eb] = 8'hca;
s_mem_contents[14'h04ec] = 8'hca;
s_mem_contents[14'h04ed] = 8'hca;
s_mem_contents[14'h04ee] = 8'hca;
s_mem_contents[14'h04ef] = 8'hca;
s_mem_contents[14'h04f0] = 8'hca;
s_mem_contents[14'h04f1] = 8'hca;
s_mem_contents[14'h04f2] = 8'hca;
s_mem_contents[14'h04f3] = 8'hca;
s_mem_contents[14'h04f4] = 8'hca;
s_mem_contents[14'h04f5] = 8'hca;
s_mem_contents[14'h04f6] = 8'hca;
s_mem_contents[14'h04f7] = 8'hca;
s_mem_contents[14'h04f8] = 8'hca;
s_mem_contents[14'h04f9] = 8'hca;
s_mem_contents[14'h04fa] = 8'hca;
s_mem_contents[14'h04fb] = 8'hca;
s_mem_contents[14'h04fc] = 8'hca;
s_mem_contents[14'h04fd] = 8'hca;
s_mem_contents[14'h04fe] = 8'hca;
s_mem_contents[14'h04ff] = 8'hca;
s_mem_contents[14'h0500] = 8'hca;
s_mem_contents[14'h0501] = 8'hca;
s_mem_contents[14'h0502] = 8'hca;
s_mem_contents[14'h0503] = 8'hca;
s_mem_contents[14'h0504] = 8'hca;
s_mem_contents[14'h0505] = 8'hca;
s_mem_contents[14'h0506] = 8'hca;
s_mem_contents[14'h0507] = 8'hca;
s_mem_contents[14'h0508] = 8'hca;
s_mem_contents[14'h0509] = 8'hca;
s_mem_contents[14'h050a] = 8'hca;
s_mem_contents[14'h050b] = 8'hca;
s_mem_contents[14'h050c] = 8'hca;
s_mem_contents[14'h050d] = 8'hca;
s_mem_contents[14'h050e] = 8'hca;
s_mem_contents[14'h050f] = 8'hca;
s_mem_contents[14'h0510] = 8'hca;
s_mem_contents[14'h0511] = 8'hca;
s_mem_contents[14'h0512] = 8'hca;
s_mem_contents[14'h0513] = 8'hca;
s_mem_contents[14'h0514] = 8'hca;
s_mem_contents[14'h0515] = 8'hca;
s_mem_contents[14'h0516] = 8'hca;
s_mem_contents[14'h0517] = 8'hca;
s_mem_contents[14'h0518] = 8'hca;
s_mem_contents[14'h0519] = 8'hca;
s_mem_contents[14'h051a] = 8'hca;
s_mem_contents[14'h051b] = 8'hca;
s_mem_contents[14'h051c] = 8'hca;
s_mem_contents[14'h051d] = 8'hca;
s_mem_contents[14'h051e] = 8'hca;
s_mem_contents[14'h051f] = 8'hca;
s_mem_contents[14'h0520] = 8'hca;
s_mem_contents[14'h0521] = 8'hca;
s_mem_contents[14'h0522] = 8'hca;
s_mem_contents[14'h0523] = 8'hca;
s_mem_contents[14'h0524] = 8'hca;
s_mem_contents[14'h0525] = 8'hca;
s_mem_contents[14'h0526] = 8'hca;
s_mem_contents[14'h0527] = 8'hca;
s_mem_contents[14'h0528] = 8'hca;
s_mem_contents[14'h0529] = 8'hca;
s_mem_contents[14'h052a] = 8'hca;
s_mem_contents[14'h052b] = 8'hca;
s_mem_contents[14'h052c] = 8'hca;
s_mem_contents[14'h052d] = 8'hca;
s_mem_contents[14'h052e] = 8'hca;
s_mem_contents[14'h052f] = 8'hca;
s_mem_contents[14'h0530] = 8'hca;
s_mem_contents[14'h0531] = 8'hca;
s_mem_contents[14'h0532] = 8'hca;
s_mem_contents[14'h0533] = 8'hca;
s_mem_contents[14'h0534] = 8'hca;
s_mem_contents[14'h0535] = 8'hca;
s_mem_contents[14'h0536] = 8'hca;
s_mem_contents[14'h0537] = 8'hca;
s_mem_contents[14'h0538] = 8'hca;
s_mem_contents[14'h0539] = 8'hca;
s_mem_contents[14'h053a] = 8'hca;
s_mem_contents[14'h053b] = 8'hca;
s_mem_contents[14'h053c] = 8'hca;
s_mem_contents[14'h053d] = 8'hca;
s_mem_contents[14'h053e] = 8'hca;
s_mem_contents[14'h053f] = 8'hca;
s_mem_contents[14'h0540] = 8'hca;
s_mem_contents[14'h0541] = 8'hca;
s_mem_contents[14'h0542] = 8'hca;
s_mem_contents[14'h0543] = 8'hca;
s_mem_contents[14'h0544] = 8'hca;
s_mem_contents[14'h0545] = 8'hca;
s_mem_contents[14'h0546] = 8'hca;
s_mem_contents[14'h0547] = 8'hca;
s_mem_contents[14'h0548] = 8'hca;
s_mem_contents[14'h0549] = 8'hca;
s_mem_contents[14'h054a] = 8'hca;
s_mem_contents[14'h054b] = 8'hca;
s_mem_contents[14'h054c] = 8'hca;
s_mem_contents[14'h054d] = 8'hca;
s_mem_contents[14'h054e] = 8'hca;
s_mem_contents[14'h054f] = 8'hca;
s_mem_contents[14'h0550] = 8'hca;
s_mem_contents[14'h0551] = 8'hca;
s_mem_contents[14'h0552] = 8'hca;
s_mem_contents[14'h0553] = 8'hca;
s_mem_contents[14'h0554] = 8'hca;
s_mem_contents[14'h0555] = 8'hca;
s_mem_contents[14'h0556] = 8'hca;
s_mem_contents[14'h0557] = 8'hca;
s_mem_contents[14'h0558] = 8'hca;
s_mem_contents[14'h0559] = 8'hca;
s_mem_contents[14'h055a] = 8'hca;
s_mem_contents[14'h055b] = 8'hca;
s_mem_contents[14'h055c] = 8'hca;
s_mem_contents[14'h055d] = 8'hca;
s_mem_contents[14'h055e] = 8'hca;
s_mem_contents[14'h055f] = 8'hca;
s_mem_contents[14'h0560] = 8'hca;
s_mem_contents[14'h0561] = 8'hca;
s_mem_contents[14'h0562] = 8'hca;
s_mem_contents[14'h0563] = 8'hca;
s_mem_contents[14'h0564] = 8'hca;
s_mem_contents[14'h0565] = 8'hca;
s_mem_contents[14'h0566] = 8'hea;
s_mem_contents[14'h0567] = 8'hea;
s_mem_contents[14'h0568] = 8'hea;
s_mem_contents[14'h0569] = 8'hea;
s_mem_contents[14'h056a] = 8'hea;
s_mem_contents[14'h056b] = 8'hf0;
s_mem_contents[14'h056c] = 8'h08;
s_mem_contents[14'h056d] = 8'h4c;
s_mem_contents[14'h056e] = 8'h6d;
s_mem_contents[14'h056f] = 8'h05;
s_mem_contents[14'h0570] = 8'hea;
s_mem_contents[14'h0571] = 8'hea;
s_mem_contents[14'h0572] = 8'hea;
s_mem_contents[14'h0573] = 8'hea;
s_mem_contents[14'h0574] = 8'hea;
s_mem_contents[14'h0575] = 8'hea;
s_mem_contents[14'h0576] = 8'hea;
s_mem_contents[14'h0577] = 8'hea;
s_mem_contents[14'h0578] = 8'hea;
s_mem_contents[14'h0579] = 8'hea;
s_mem_contents[14'h057a] = 8'hc0;
s_mem_contents[14'h057b] = 8'h00;
s_mem_contents[14'h057c] = 8'hf0;
s_mem_contents[14'h057d] = 8'h03;
s_mem_contents[14'h057e] = 8'h4c;
s_mem_contents[14'h057f] = 8'h46;
s_mem_contents[14'h0580] = 8'h04;
s_mem_contents[14'h0581] = 8'had;
s_mem_contents[14'h0582] = 8'h00;
s_mem_contents[14'h0583] = 8'h02;
s_mem_contents[14'h0584] = 8'hc9;
s_mem_contents[14'h0585] = 8'h01;
s_mem_contents[14'h0586] = 8'hd0;
s_mem_contents[14'h0587] = 8'hfe;
s_mem_contents[14'h0588] = 8'ha9;
s_mem_contents[14'h0589] = 8'h02;
s_mem_contents[14'h058a] = 8'h8d;
s_mem_contents[14'h058b] = 8'h00;
s_mem_contents[14'h058c] = 8'h02;
s_mem_contents[14'h058d] = 8'hc0;
s_mem_contents[14'h058e] = 8'h01;
s_mem_contents[14'h058f] = 8'hd0;
s_mem_contents[14'h0590] = 8'h03;
s_mem_contents[14'h0591] = 8'h4c;
s_mem_contents[14'h0592] = 8'h91;
s_mem_contents[14'h0593] = 8'h05;
s_mem_contents[14'h0594] = 8'ha9;
s_mem_contents[14'h0595] = 8'h00;
s_mem_contents[14'h0596] = 8'hc9;
s_mem_contents[14'h0597] = 8'h00;
s_mem_contents[14'h0598] = 8'hd0;
s_mem_contents[14'h0599] = 8'hfe;
s_mem_contents[14'h059a] = 8'h90;
s_mem_contents[14'h059b] = 8'hfe;
s_mem_contents[14'h059c] = 8'h30;
s_mem_contents[14'h059d] = 8'hfe;
s_mem_contents[14'h059e] = 8'hc9;
s_mem_contents[14'h059f] = 8'h01;
s_mem_contents[14'h05a0] = 8'hf0;
s_mem_contents[14'h05a1] = 8'hfe;
s_mem_contents[14'h05a2] = 8'hb0;
s_mem_contents[14'h05a3] = 8'hfe;
s_mem_contents[14'h05a4] = 8'h10;
s_mem_contents[14'h05a5] = 8'hfe;
s_mem_contents[14'h05a6] = 8'haa;
s_mem_contents[14'h05a7] = 8'he0;
s_mem_contents[14'h05a8] = 8'h00;
s_mem_contents[14'h05a9] = 8'hd0;
s_mem_contents[14'h05aa] = 8'hfe;
s_mem_contents[14'h05ab] = 8'h90;
s_mem_contents[14'h05ac] = 8'hfe;
s_mem_contents[14'h05ad] = 8'h30;
s_mem_contents[14'h05ae] = 8'hfe;
s_mem_contents[14'h05af] = 8'he0;
s_mem_contents[14'h05b0] = 8'h01;
s_mem_contents[14'h05b1] = 8'hf0;
s_mem_contents[14'h05b2] = 8'hfe;
s_mem_contents[14'h05b3] = 8'hb0;
s_mem_contents[14'h05b4] = 8'hfe;
s_mem_contents[14'h05b5] = 8'h10;
s_mem_contents[14'h05b6] = 8'hfe;
s_mem_contents[14'h05b7] = 8'ha8;
s_mem_contents[14'h05b8] = 8'hc0;
s_mem_contents[14'h05b9] = 8'h00;
s_mem_contents[14'h05ba] = 8'hd0;
s_mem_contents[14'h05bb] = 8'hfe;
s_mem_contents[14'h05bc] = 8'h90;
s_mem_contents[14'h05bd] = 8'hfe;
s_mem_contents[14'h05be] = 8'h30;
s_mem_contents[14'h05bf] = 8'hfe;
s_mem_contents[14'h05c0] = 8'hc0;
s_mem_contents[14'h05c1] = 8'h01;
s_mem_contents[14'h05c2] = 8'hf0;
s_mem_contents[14'h05c3] = 8'hfe;
s_mem_contents[14'h05c4] = 8'hb0;
s_mem_contents[14'h05c5] = 8'hfe;
s_mem_contents[14'h05c6] = 8'h10;
s_mem_contents[14'h05c7] = 8'hfe;
s_mem_contents[14'h05c8] = 8'had;
s_mem_contents[14'h05c9] = 8'h00;
s_mem_contents[14'h05ca] = 8'h02;
s_mem_contents[14'h05cb] = 8'hc9;
s_mem_contents[14'h05cc] = 8'h02;
s_mem_contents[14'h05cd] = 8'hd0;
s_mem_contents[14'h05ce] = 8'hfe;
s_mem_contents[14'h05cf] = 8'ha9;
s_mem_contents[14'h05d0] = 8'h03;
s_mem_contents[14'h05d1] = 8'h8d;
s_mem_contents[14'h05d2] = 8'h00;
s_mem_contents[14'h05d3] = 8'h02;
s_mem_contents[14'h05d4] = 8'ha2;
s_mem_contents[14'h05d5] = 8'hff;
s_mem_contents[14'h05d6] = 8'h9a;
s_mem_contents[14'h05d7] = 8'ha9;
s_mem_contents[14'h05d8] = 8'h55;
s_mem_contents[14'h05d9] = 8'h48;
s_mem_contents[14'h05da] = 8'ha9;
s_mem_contents[14'h05db] = 8'haa;
s_mem_contents[14'h05dc] = 8'h48;
s_mem_contents[14'h05dd] = 8'hcd;
s_mem_contents[14'h05de] = 8'hfe;
s_mem_contents[14'h05df] = 8'h01;
s_mem_contents[14'h05e0] = 8'hd0;
s_mem_contents[14'h05e1] = 8'hfe;
s_mem_contents[14'h05e2] = 8'hba;
s_mem_contents[14'h05e3] = 8'h8a;
s_mem_contents[14'h05e4] = 8'hc9;
s_mem_contents[14'h05e5] = 8'hfd;
s_mem_contents[14'h05e6] = 8'hd0;
s_mem_contents[14'h05e7] = 8'hfe;
s_mem_contents[14'h05e8] = 8'h68;
s_mem_contents[14'h05e9] = 8'hc9;
s_mem_contents[14'h05ea] = 8'haa;
s_mem_contents[14'h05eb] = 8'hd0;
s_mem_contents[14'h05ec] = 8'hfe;
s_mem_contents[14'h05ed] = 8'h68;
s_mem_contents[14'h05ee] = 8'hc9;
s_mem_contents[14'h05ef] = 8'h55;
s_mem_contents[14'h05f0] = 8'hd0;
s_mem_contents[14'h05f1] = 8'hfe;
s_mem_contents[14'h05f2] = 8'hcd;
s_mem_contents[14'h05f3] = 8'hff;
s_mem_contents[14'h05f4] = 8'h01;
s_mem_contents[14'h05f5] = 8'hd0;
s_mem_contents[14'h05f6] = 8'hfe;
s_mem_contents[14'h05f7] = 8'hba;
s_mem_contents[14'h05f8] = 8'he0;
s_mem_contents[14'h05f9] = 8'hff;
s_mem_contents[14'h05fa] = 8'hd0;
s_mem_contents[14'h05fb] = 8'hfe;
s_mem_contents[14'h05fc] = 8'had;
s_mem_contents[14'h05fd] = 8'h00;
s_mem_contents[14'h05fe] = 8'h02;
s_mem_contents[14'h05ff] = 8'hc9;
s_mem_contents[14'h0600] = 8'h03;
s_mem_contents[14'h0601] = 8'hd0;
s_mem_contents[14'h0602] = 8'hfe;
s_mem_contents[14'h0603] = 8'ha9;
s_mem_contents[14'h0604] = 8'h04;
s_mem_contents[14'h0605] = 8'h8d;
s_mem_contents[14'h0606] = 8'h00;
s_mem_contents[14'h0607] = 8'h02;
s_mem_contents[14'h0608] = 8'ha9;
s_mem_contents[14'h0609] = 8'hff;
s_mem_contents[14'h060a] = 8'h48;
s_mem_contents[14'h060b] = 8'h28;
s_mem_contents[14'h060c] = 8'h10;
s_mem_contents[14'h060d] = 8'h1a;
s_mem_contents[14'h060e] = 8'h50;
s_mem_contents[14'h060f] = 8'h1b;
s_mem_contents[14'h0610] = 8'h90;
s_mem_contents[14'h0611] = 8'h1c;
s_mem_contents[14'h0612] = 8'hd0;
s_mem_contents[14'h0613] = 8'h1d;
s_mem_contents[14'h0614] = 8'h30;
s_mem_contents[14'h0615] = 8'h03;
s_mem_contents[14'h0616] = 8'h4c;
s_mem_contents[14'h0617] = 8'h16;
s_mem_contents[14'h0618] = 8'h06;
s_mem_contents[14'h0619] = 8'h70;
s_mem_contents[14'h061a] = 8'h03;
s_mem_contents[14'h061b] = 8'h4c;
s_mem_contents[14'h061c] = 8'h1b;
s_mem_contents[14'h061d] = 8'h06;
s_mem_contents[14'h061e] = 8'hb0;
s_mem_contents[14'h061f] = 8'h03;
s_mem_contents[14'h0620] = 8'h4c;
s_mem_contents[14'h0621] = 8'h20;
s_mem_contents[14'h0622] = 8'h06;
s_mem_contents[14'h0623] = 8'hf0;
s_mem_contents[14'h0624] = 8'h0f;
s_mem_contents[14'h0625] = 8'h4c;
s_mem_contents[14'h0626] = 8'h25;
s_mem_contents[14'h0627] = 8'h06;
s_mem_contents[14'h0628] = 8'h4c;
s_mem_contents[14'h0629] = 8'h28;
s_mem_contents[14'h062a] = 8'h06;
s_mem_contents[14'h062b] = 8'h4c;
s_mem_contents[14'h062c] = 8'h2b;
s_mem_contents[14'h062d] = 8'h06;
s_mem_contents[14'h062e] = 8'h4c;
s_mem_contents[14'h062f] = 8'h2e;
s_mem_contents[14'h0630] = 8'h06;
s_mem_contents[14'h0631] = 8'h4c;
s_mem_contents[14'h0632] = 8'h31;
s_mem_contents[14'h0633] = 8'h06;
s_mem_contents[14'h0634] = 8'h08;
s_mem_contents[14'h0635] = 8'hba;
s_mem_contents[14'h0636] = 8'he0;
s_mem_contents[14'h0637] = 8'hfe;
s_mem_contents[14'h0638] = 8'hd0;
s_mem_contents[14'h0639] = 8'hfe;
s_mem_contents[14'h063a] = 8'h68;
s_mem_contents[14'h063b] = 8'hc9;
s_mem_contents[14'h063c] = 8'hff;
s_mem_contents[14'h063d] = 8'hd0;
s_mem_contents[14'h063e] = 8'hfe;
s_mem_contents[14'h063f] = 8'hba;
s_mem_contents[14'h0640] = 8'he0;
s_mem_contents[14'h0641] = 8'hff;
s_mem_contents[14'h0642] = 8'hd0;
s_mem_contents[14'h0643] = 8'hfe;
s_mem_contents[14'h0644] = 8'ha9;
s_mem_contents[14'h0645] = 8'h00;
s_mem_contents[14'h0646] = 8'h48;
s_mem_contents[14'h0647] = 8'h28;
s_mem_contents[14'h0648] = 8'h30;
s_mem_contents[14'h0649] = 8'h1a;
s_mem_contents[14'h064a] = 8'h70;
s_mem_contents[14'h064b] = 8'h1b;
s_mem_contents[14'h064c] = 8'hb0;
s_mem_contents[14'h064d] = 8'h1c;
s_mem_contents[14'h064e] = 8'hf0;
s_mem_contents[14'h064f] = 8'h1d;
s_mem_contents[14'h0650] = 8'h10;
s_mem_contents[14'h0651] = 8'h03;
s_mem_contents[14'h0652] = 8'h4c;
s_mem_contents[14'h0653] = 8'h52;
s_mem_contents[14'h0654] = 8'h06;
s_mem_contents[14'h0655] = 8'h50;
s_mem_contents[14'h0656] = 8'h03;
s_mem_contents[14'h0657] = 8'h4c;
s_mem_contents[14'h0658] = 8'h57;
s_mem_contents[14'h0659] = 8'h06;
s_mem_contents[14'h065a] = 8'h90;
s_mem_contents[14'h065b] = 8'h03;
s_mem_contents[14'h065c] = 8'h4c;
s_mem_contents[14'h065d] = 8'h5c;
s_mem_contents[14'h065e] = 8'h06;
s_mem_contents[14'h065f] = 8'hd0;
s_mem_contents[14'h0660] = 8'h0f;
s_mem_contents[14'h0661] = 8'h4c;
s_mem_contents[14'h0662] = 8'h61;
s_mem_contents[14'h0663] = 8'h06;
s_mem_contents[14'h0664] = 8'h4c;
s_mem_contents[14'h0665] = 8'h64;
s_mem_contents[14'h0666] = 8'h06;
s_mem_contents[14'h0667] = 8'h4c;
s_mem_contents[14'h0668] = 8'h67;
s_mem_contents[14'h0669] = 8'h06;
s_mem_contents[14'h066a] = 8'h4c;
s_mem_contents[14'h066b] = 8'h6a;
s_mem_contents[14'h066c] = 8'h06;
s_mem_contents[14'h066d] = 8'h4c;
s_mem_contents[14'h066e] = 8'h6d;
s_mem_contents[14'h066f] = 8'h06;
s_mem_contents[14'h0670] = 8'h08;
s_mem_contents[14'h0671] = 8'h68;
s_mem_contents[14'h0672] = 8'hc9;
s_mem_contents[14'h0673] = 8'h30;
s_mem_contents[14'h0674] = 8'hd0;
s_mem_contents[14'h0675] = 8'hfe;
s_mem_contents[14'h0676] = 8'ha9;
s_mem_contents[14'h0677] = 8'h02;
s_mem_contents[14'h0678] = 8'h48;
s_mem_contents[14'h0679] = 8'h28;
s_mem_contents[14'h067a] = 8'hd0;
s_mem_contents[14'h067b] = 8'h02;
s_mem_contents[14'h067c] = 8'hf0;
s_mem_contents[14'h067d] = 8'h03;
s_mem_contents[14'h067e] = 8'h4c;
s_mem_contents[14'h067f] = 8'h7e;
s_mem_contents[14'h0680] = 8'h06;
s_mem_contents[14'h0681] = 8'hb0;
s_mem_contents[14'h0682] = 8'h02;
s_mem_contents[14'h0683] = 8'h90;
s_mem_contents[14'h0684] = 8'h03;
s_mem_contents[14'h0685] = 8'h4c;
s_mem_contents[14'h0686] = 8'h85;
s_mem_contents[14'h0687] = 8'h06;
s_mem_contents[14'h0688] = 8'h30;
s_mem_contents[14'h0689] = 8'h02;
s_mem_contents[14'h068a] = 8'h10;
s_mem_contents[14'h068b] = 8'h03;
s_mem_contents[14'h068c] = 8'h4c;
s_mem_contents[14'h068d] = 8'h8c;
s_mem_contents[14'h068e] = 8'h06;
s_mem_contents[14'h068f] = 8'h70;
s_mem_contents[14'h0690] = 8'h02;
s_mem_contents[14'h0691] = 8'h50;
s_mem_contents[14'h0692] = 8'h03;
s_mem_contents[14'h0693] = 8'h4c;
s_mem_contents[14'h0694] = 8'h93;
s_mem_contents[14'h0695] = 8'h06;
s_mem_contents[14'h0696] = 8'ha9;
s_mem_contents[14'h0697] = 8'h01;
s_mem_contents[14'h0698] = 8'h48;
s_mem_contents[14'h0699] = 8'h28;
s_mem_contents[14'h069a] = 8'hf0;
s_mem_contents[14'h069b] = 8'h02;
s_mem_contents[14'h069c] = 8'hd0;
s_mem_contents[14'h069d] = 8'h03;
s_mem_contents[14'h069e] = 8'h4c;
s_mem_contents[14'h069f] = 8'h9e;
s_mem_contents[14'h06a0] = 8'h06;
s_mem_contents[14'h06a1] = 8'h90;
s_mem_contents[14'h06a2] = 8'h02;
s_mem_contents[14'h06a3] = 8'hb0;
s_mem_contents[14'h06a4] = 8'h03;
s_mem_contents[14'h06a5] = 8'h4c;
s_mem_contents[14'h06a6] = 8'ha5;
s_mem_contents[14'h06a7] = 8'h06;
s_mem_contents[14'h06a8] = 8'h30;
s_mem_contents[14'h06a9] = 8'h02;
s_mem_contents[14'h06aa] = 8'h10;
s_mem_contents[14'h06ab] = 8'h03;
s_mem_contents[14'h06ac] = 8'h4c;
s_mem_contents[14'h06ad] = 8'hac;
s_mem_contents[14'h06ae] = 8'h06;
s_mem_contents[14'h06af] = 8'h70;
s_mem_contents[14'h06b0] = 8'h02;
s_mem_contents[14'h06b1] = 8'h50;
s_mem_contents[14'h06b2] = 8'h03;
s_mem_contents[14'h06b3] = 8'h4c;
s_mem_contents[14'h06b4] = 8'hb3;
s_mem_contents[14'h06b5] = 8'h06;
s_mem_contents[14'h06b6] = 8'ha9;
s_mem_contents[14'h06b7] = 8'h80;
s_mem_contents[14'h06b8] = 8'h48;
s_mem_contents[14'h06b9] = 8'h28;
s_mem_contents[14'h06ba] = 8'hf0;
s_mem_contents[14'h06bb] = 8'h02;
s_mem_contents[14'h06bc] = 8'hd0;
s_mem_contents[14'h06bd] = 8'h03;
s_mem_contents[14'h06be] = 8'h4c;
s_mem_contents[14'h06bf] = 8'hbe;
s_mem_contents[14'h06c0] = 8'h06;
s_mem_contents[14'h06c1] = 8'hb0;
s_mem_contents[14'h06c2] = 8'h02;
s_mem_contents[14'h06c3] = 8'h90;
s_mem_contents[14'h06c4] = 8'h03;
s_mem_contents[14'h06c5] = 8'h4c;
s_mem_contents[14'h06c6] = 8'hc5;
s_mem_contents[14'h06c7] = 8'h06;
s_mem_contents[14'h06c8] = 8'h10;
s_mem_contents[14'h06c9] = 8'h02;
s_mem_contents[14'h06ca] = 8'h30;
s_mem_contents[14'h06cb] = 8'h03;
s_mem_contents[14'h06cc] = 8'h4c;
s_mem_contents[14'h06cd] = 8'hcc;
s_mem_contents[14'h06ce] = 8'h06;
s_mem_contents[14'h06cf] = 8'h70;
s_mem_contents[14'h06d0] = 8'h02;
s_mem_contents[14'h06d1] = 8'h50;
s_mem_contents[14'h06d2] = 8'h03;
s_mem_contents[14'h06d3] = 8'h4c;
s_mem_contents[14'h06d4] = 8'hd3;
s_mem_contents[14'h06d5] = 8'h06;
s_mem_contents[14'h06d6] = 8'ha9;
s_mem_contents[14'h06d7] = 8'h40;
s_mem_contents[14'h06d8] = 8'h48;
s_mem_contents[14'h06d9] = 8'h28;
s_mem_contents[14'h06da] = 8'hf0;
s_mem_contents[14'h06db] = 8'h02;
s_mem_contents[14'h06dc] = 8'hd0;
s_mem_contents[14'h06dd] = 8'h03;
s_mem_contents[14'h06de] = 8'h4c;
s_mem_contents[14'h06df] = 8'hde;
s_mem_contents[14'h06e0] = 8'h06;
s_mem_contents[14'h06e1] = 8'hb0;
s_mem_contents[14'h06e2] = 8'h02;
s_mem_contents[14'h06e3] = 8'h90;
s_mem_contents[14'h06e4] = 8'h03;
s_mem_contents[14'h06e5] = 8'h4c;
s_mem_contents[14'h06e6] = 8'he5;
s_mem_contents[14'h06e7] = 8'h06;
s_mem_contents[14'h06e8] = 8'h30;
s_mem_contents[14'h06e9] = 8'h02;
s_mem_contents[14'h06ea] = 8'h10;
s_mem_contents[14'h06eb] = 8'h03;
s_mem_contents[14'h06ec] = 8'h4c;
s_mem_contents[14'h06ed] = 8'hec;
s_mem_contents[14'h06ee] = 8'h06;
s_mem_contents[14'h06ef] = 8'h50;
s_mem_contents[14'h06f0] = 8'h02;
s_mem_contents[14'h06f1] = 8'h70;
s_mem_contents[14'h06f2] = 8'h03;
s_mem_contents[14'h06f3] = 8'h4c;
s_mem_contents[14'h06f4] = 8'hf3;
s_mem_contents[14'h06f5] = 8'h06;
s_mem_contents[14'h06f6] = 8'ha9;
s_mem_contents[14'h06f7] = 8'hfd;
s_mem_contents[14'h06f8] = 8'h48;
s_mem_contents[14'h06f9] = 8'h28;
s_mem_contents[14'h06fa] = 8'hf0;
s_mem_contents[14'h06fb] = 8'h02;
s_mem_contents[14'h06fc] = 8'hd0;
s_mem_contents[14'h06fd] = 8'h03;
s_mem_contents[14'h06fe] = 8'h4c;
s_mem_contents[14'h06ff] = 8'hfe;
s_mem_contents[14'h0700] = 8'h06;
s_mem_contents[14'h0701] = 8'h90;
s_mem_contents[14'h0702] = 8'h02;
s_mem_contents[14'h0703] = 8'hb0;
s_mem_contents[14'h0704] = 8'h03;
s_mem_contents[14'h0705] = 8'h4c;
s_mem_contents[14'h0706] = 8'h05;
s_mem_contents[14'h0707] = 8'h07;
s_mem_contents[14'h0708] = 8'h10;
s_mem_contents[14'h0709] = 8'h02;
s_mem_contents[14'h070a] = 8'h30;
s_mem_contents[14'h070b] = 8'h03;
s_mem_contents[14'h070c] = 8'h4c;
s_mem_contents[14'h070d] = 8'h0c;
s_mem_contents[14'h070e] = 8'h07;
s_mem_contents[14'h070f] = 8'h50;
s_mem_contents[14'h0710] = 8'h02;
s_mem_contents[14'h0711] = 8'h70;
s_mem_contents[14'h0712] = 8'h03;
s_mem_contents[14'h0713] = 8'h4c;
s_mem_contents[14'h0714] = 8'h13;
s_mem_contents[14'h0715] = 8'h07;
s_mem_contents[14'h0716] = 8'ha9;
s_mem_contents[14'h0717] = 8'hfe;
s_mem_contents[14'h0718] = 8'h48;
s_mem_contents[14'h0719] = 8'h28;
s_mem_contents[14'h071a] = 8'hd0;
s_mem_contents[14'h071b] = 8'h02;
s_mem_contents[14'h071c] = 8'hf0;
s_mem_contents[14'h071d] = 8'h03;
s_mem_contents[14'h071e] = 8'h4c;
s_mem_contents[14'h071f] = 8'h1e;
s_mem_contents[14'h0720] = 8'h07;
s_mem_contents[14'h0721] = 8'hb0;
s_mem_contents[14'h0722] = 8'h02;
s_mem_contents[14'h0723] = 8'h90;
s_mem_contents[14'h0724] = 8'h03;
s_mem_contents[14'h0725] = 8'h4c;
s_mem_contents[14'h0726] = 8'h25;
s_mem_contents[14'h0727] = 8'h07;
s_mem_contents[14'h0728] = 8'h10;
s_mem_contents[14'h0729] = 8'h02;
s_mem_contents[14'h072a] = 8'h30;
s_mem_contents[14'h072b] = 8'h03;
s_mem_contents[14'h072c] = 8'h4c;
s_mem_contents[14'h072d] = 8'h2c;
s_mem_contents[14'h072e] = 8'h07;
s_mem_contents[14'h072f] = 8'h50;
s_mem_contents[14'h0730] = 8'h02;
s_mem_contents[14'h0731] = 8'h70;
s_mem_contents[14'h0732] = 8'h03;
s_mem_contents[14'h0733] = 8'h4c;
s_mem_contents[14'h0734] = 8'h33;
s_mem_contents[14'h0735] = 8'h07;
s_mem_contents[14'h0736] = 8'ha9;
s_mem_contents[14'h0737] = 8'h7f;
s_mem_contents[14'h0738] = 8'h48;
s_mem_contents[14'h0739] = 8'h28;
s_mem_contents[14'h073a] = 8'hd0;
s_mem_contents[14'h073b] = 8'h02;
s_mem_contents[14'h073c] = 8'hf0;
s_mem_contents[14'h073d] = 8'h03;
s_mem_contents[14'h073e] = 8'h4c;
s_mem_contents[14'h073f] = 8'h3e;
s_mem_contents[14'h0740] = 8'h07;
s_mem_contents[14'h0741] = 8'h90;
s_mem_contents[14'h0742] = 8'h02;
s_mem_contents[14'h0743] = 8'hb0;
s_mem_contents[14'h0744] = 8'h03;
s_mem_contents[14'h0745] = 8'h4c;
s_mem_contents[14'h0746] = 8'h45;
s_mem_contents[14'h0747] = 8'h07;
s_mem_contents[14'h0748] = 8'h30;
s_mem_contents[14'h0749] = 8'h02;
s_mem_contents[14'h074a] = 8'h10;
s_mem_contents[14'h074b] = 8'h03;
s_mem_contents[14'h074c] = 8'h4c;
s_mem_contents[14'h074d] = 8'h4c;
s_mem_contents[14'h074e] = 8'h07;
s_mem_contents[14'h074f] = 8'h50;
s_mem_contents[14'h0750] = 8'h02;
s_mem_contents[14'h0751] = 8'h70;
s_mem_contents[14'h0752] = 8'h03;
s_mem_contents[14'h0753] = 8'h4c;
s_mem_contents[14'h0754] = 8'h53;
s_mem_contents[14'h0755] = 8'h07;
s_mem_contents[14'h0756] = 8'ha9;
s_mem_contents[14'h0757] = 8'hbf;
s_mem_contents[14'h0758] = 8'h48;
s_mem_contents[14'h0759] = 8'h28;
s_mem_contents[14'h075a] = 8'hd0;
s_mem_contents[14'h075b] = 8'h02;
s_mem_contents[14'h075c] = 8'hf0;
s_mem_contents[14'h075d] = 8'h03;
s_mem_contents[14'h075e] = 8'h4c;
s_mem_contents[14'h075f] = 8'h5e;
s_mem_contents[14'h0760] = 8'h07;
s_mem_contents[14'h0761] = 8'h90;
s_mem_contents[14'h0762] = 8'h02;
s_mem_contents[14'h0763] = 8'hb0;
s_mem_contents[14'h0764] = 8'h03;
s_mem_contents[14'h0765] = 8'h4c;
s_mem_contents[14'h0766] = 8'h65;
s_mem_contents[14'h0767] = 8'h07;
s_mem_contents[14'h0768] = 8'h10;
s_mem_contents[14'h0769] = 8'h02;
s_mem_contents[14'h076a] = 8'h30;
s_mem_contents[14'h076b] = 8'h03;
s_mem_contents[14'h076c] = 8'h4c;
s_mem_contents[14'h076d] = 8'h6c;
s_mem_contents[14'h076e] = 8'h07;
s_mem_contents[14'h076f] = 8'h70;
s_mem_contents[14'h0770] = 8'h02;
s_mem_contents[14'h0771] = 8'h50;
s_mem_contents[14'h0772] = 8'h03;
s_mem_contents[14'h0773] = 8'h4c;
s_mem_contents[14'h0774] = 8'h73;
s_mem_contents[14'h0775] = 8'h07;
s_mem_contents[14'h0776] = 8'had;
s_mem_contents[14'h0777] = 8'h00;
s_mem_contents[14'h0778] = 8'h02;
s_mem_contents[14'h0779] = 8'hc9;
s_mem_contents[14'h077a] = 8'h04;
s_mem_contents[14'h077b] = 8'hd0;
s_mem_contents[14'h077c] = 8'hfe;
s_mem_contents[14'h077d] = 8'ha9;
s_mem_contents[14'h077e] = 8'h05;
s_mem_contents[14'h077f] = 8'h8d;
s_mem_contents[14'h0780] = 8'h00;
s_mem_contents[14'h0781] = 8'h02;
s_mem_contents[14'h0782] = 8'ha2;
s_mem_contents[14'h0783] = 8'h55;
s_mem_contents[14'h0784] = 8'ha0;
s_mem_contents[14'h0785] = 8'haa;
s_mem_contents[14'h0786] = 8'ha9;
s_mem_contents[14'h0787] = 8'hff;
s_mem_contents[14'h0788] = 8'h48;
s_mem_contents[14'h0789] = 8'ha9;
s_mem_contents[14'h078a] = 8'h01;
s_mem_contents[14'h078b] = 8'h28;
s_mem_contents[14'h078c] = 8'h48;
s_mem_contents[14'h078d] = 8'h08;
s_mem_contents[14'h078e] = 8'hc9;
s_mem_contents[14'h078f] = 8'h01;
s_mem_contents[14'h0790] = 8'hd0;
s_mem_contents[14'h0791] = 8'hfe;
s_mem_contents[14'h0792] = 8'h68;
s_mem_contents[14'h0793] = 8'h48;
s_mem_contents[14'h0794] = 8'hc9;
s_mem_contents[14'h0795] = 8'hff;
s_mem_contents[14'h0796] = 8'hd0;
s_mem_contents[14'h0797] = 8'hfe;
s_mem_contents[14'h0798] = 8'h28;
s_mem_contents[14'h0799] = 8'ha9;
s_mem_contents[14'h079a] = 8'h00;
s_mem_contents[14'h079b] = 8'h48;
s_mem_contents[14'h079c] = 8'ha9;
s_mem_contents[14'h079d] = 8'h00;
s_mem_contents[14'h079e] = 8'h28;
s_mem_contents[14'h079f] = 8'h48;
s_mem_contents[14'h07a0] = 8'h08;
s_mem_contents[14'h07a1] = 8'hc9;
s_mem_contents[14'h07a2] = 8'h00;
s_mem_contents[14'h07a3] = 8'hd0;
s_mem_contents[14'h07a4] = 8'hfe;
s_mem_contents[14'h07a5] = 8'h68;
s_mem_contents[14'h07a6] = 8'h48;
s_mem_contents[14'h07a7] = 8'hc9;
s_mem_contents[14'h07a8] = 8'h30;
s_mem_contents[14'h07a9] = 8'hd0;
s_mem_contents[14'h07aa] = 8'hfe;
s_mem_contents[14'h07ab] = 8'h28;
s_mem_contents[14'h07ac] = 8'ha9;
s_mem_contents[14'h07ad] = 8'hff;
s_mem_contents[14'h07ae] = 8'h48;
s_mem_contents[14'h07af] = 8'ha9;
s_mem_contents[14'h07b0] = 8'hff;
s_mem_contents[14'h07b1] = 8'h28;
s_mem_contents[14'h07b2] = 8'h48;
s_mem_contents[14'h07b3] = 8'h08;
s_mem_contents[14'h07b4] = 8'hc9;
s_mem_contents[14'h07b5] = 8'hff;
s_mem_contents[14'h07b6] = 8'hd0;
s_mem_contents[14'h07b7] = 8'hfe;
s_mem_contents[14'h07b8] = 8'h68;
s_mem_contents[14'h07b9] = 8'h48;
s_mem_contents[14'h07ba] = 8'hc9;
s_mem_contents[14'h07bb] = 8'hff;
s_mem_contents[14'h07bc] = 8'hd0;
s_mem_contents[14'h07bd] = 8'hfe;
s_mem_contents[14'h07be] = 8'h28;
s_mem_contents[14'h07bf] = 8'ha9;
s_mem_contents[14'h07c0] = 8'h00;
s_mem_contents[14'h07c1] = 8'h48;
s_mem_contents[14'h07c2] = 8'ha9;
s_mem_contents[14'h07c3] = 8'h01;
s_mem_contents[14'h07c4] = 8'h28;
s_mem_contents[14'h07c5] = 8'h48;
s_mem_contents[14'h07c6] = 8'h08;
s_mem_contents[14'h07c7] = 8'hc9;
s_mem_contents[14'h07c8] = 8'h01;
s_mem_contents[14'h07c9] = 8'hd0;
s_mem_contents[14'h07ca] = 8'hfe;
s_mem_contents[14'h07cb] = 8'h68;
s_mem_contents[14'h07cc] = 8'h48;
s_mem_contents[14'h07cd] = 8'hc9;
s_mem_contents[14'h07ce] = 8'h30;
s_mem_contents[14'h07cf] = 8'hd0;
s_mem_contents[14'h07d0] = 8'hfe;
s_mem_contents[14'h07d1] = 8'h28;
s_mem_contents[14'h07d2] = 8'ha9;
s_mem_contents[14'h07d3] = 8'hff;
s_mem_contents[14'h07d4] = 8'h48;
s_mem_contents[14'h07d5] = 8'ha9;
s_mem_contents[14'h07d6] = 8'h00;
s_mem_contents[14'h07d7] = 8'h28;
s_mem_contents[14'h07d8] = 8'h48;
s_mem_contents[14'h07d9] = 8'h08;
s_mem_contents[14'h07da] = 8'hc9;
s_mem_contents[14'h07db] = 8'h00;
s_mem_contents[14'h07dc] = 8'hd0;
s_mem_contents[14'h07dd] = 8'hfe;
s_mem_contents[14'h07de] = 8'h68;
s_mem_contents[14'h07df] = 8'h48;
s_mem_contents[14'h07e0] = 8'hc9;
s_mem_contents[14'h07e1] = 8'hff;
s_mem_contents[14'h07e2] = 8'hd0;
s_mem_contents[14'h07e3] = 8'hfe;
s_mem_contents[14'h07e4] = 8'h28;
s_mem_contents[14'h07e5] = 8'ha9;
s_mem_contents[14'h07e6] = 8'h00;
s_mem_contents[14'h07e7] = 8'h48;
s_mem_contents[14'h07e8] = 8'ha9;
s_mem_contents[14'h07e9] = 8'hff;
s_mem_contents[14'h07ea] = 8'h28;
s_mem_contents[14'h07eb] = 8'h48;
s_mem_contents[14'h07ec] = 8'h08;
s_mem_contents[14'h07ed] = 8'hc9;
s_mem_contents[14'h07ee] = 8'hff;
s_mem_contents[14'h07ef] = 8'hd0;
s_mem_contents[14'h07f0] = 8'hfe;
s_mem_contents[14'h07f1] = 8'h68;
s_mem_contents[14'h07f2] = 8'h48;
s_mem_contents[14'h07f3] = 8'hc9;
s_mem_contents[14'h07f4] = 8'h30;
s_mem_contents[14'h07f5] = 8'hd0;
s_mem_contents[14'h07f6] = 8'hfe;
s_mem_contents[14'h07f7] = 8'h28;
s_mem_contents[14'h07f8] = 8'ha9;
s_mem_contents[14'h07f9] = 8'hff;
s_mem_contents[14'h07fa] = 8'h48;
s_mem_contents[14'h07fb] = 8'ha9;
s_mem_contents[14'h07fc] = 8'h00;
s_mem_contents[14'h07fd] = 8'h28;
s_mem_contents[14'h07fe] = 8'h68;
s_mem_contents[14'h07ff] = 8'h08;
s_mem_contents[14'h0800] = 8'hc9;
s_mem_contents[14'h0801] = 8'hff;
s_mem_contents[14'h0802] = 8'hd0;
s_mem_contents[14'h0803] = 8'hfe;
s_mem_contents[14'h0804] = 8'h68;
s_mem_contents[14'h0805] = 8'h48;
s_mem_contents[14'h0806] = 8'hc9;
s_mem_contents[14'h0807] = 8'hfd;
s_mem_contents[14'h0808] = 8'hd0;
s_mem_contents[14'h0809] = 8'hfe;
s_mem_contents[14'h080a] = 8'h28;
s_mem_contents[14'h080b] = 8'ha9;
s_mem_contents[14'h080c] = 8'h00;
s_mem_contents[14'h080d] = 8'h48;
s_mem_contents[14'h080e] = 8'ha9;
s_mem_contents[14'h080f] = 8'hff;
s_mem_contents[14'h0810] = 8'h28;
s_mem_contents[14'h0811] = 8'h68;
s_mem_contents[14'h0812] = 8'h08;
s_mem_contents[14'h0813] = 8'hc9;
s_mem_contents[14'h0814] = 8'h00;
s_mem_contents[14'h0815] = 8'hd0;
s_mem_contents[14'h0816] = 8'hfe;
s_mem_contents[14'h0817] = 8'h68;
s_mem_contents[14'h0818] = 8'h48;
s_mem_contents[14'h0819] = 8'hc9;
s_mem_contents[14'h081a] = 8'h32;
s_mem_contents[14'h081b] = 8'hd0;
s_mem_contents[14'h081c] = 8'hfe;
s_mem_contents[14'h081d] = 8'h28;
s_mem_contents[14'h081e] = 8'ha9;
s_mem_contents[14'h081f] = 8'hff;
s_mem_contents[14'h0820] = 8'h48;
s_mem_contents[14'h0821] = 8'ha9;
s_mem_contents[14'h0822] = 8'hfe;
s_mem_contents[14'h0823] = 8'h28;
s_mem_contents[14'h0824] = 8'h68;
s_mem_contents[14'h0825] = 8'h08;
s_mem_contents[14'h0826] = 8'hc9;
s_mem_contents[14'h0827] = 8'h01;
s_mem_contents[14'h0828] = 8'hd0;
s_mem_contents[14'h0829] = 8'hfe;
s_mem_contents[14'h082a] = 8'h68;
s_mem_contents[14'h082b] = 8'h48;
s_mem_contents[14'h082c] = 8'hc9;
s_mem_contents[14'h082d] = 8'h7d;
s_mem_contents[14'h082e] = 8'hd0;
s_mem_contents[14'h082f] = 8'hfe;
s_mem_contents[14'h0830] = 8'h28;
s_mem_contents[14'h0831] = 8'ha9;
s_mem_contents[14'h0832] = 8'h00;
s_mem_contents[14'h0833] = 8'h48;
s_mem_contents[14'h0834] = 8'ha9;
s_mem_contents[14'h0835] = 8'h00;
s_mem_contents[14'h0836] = 8'h28;
s_mem_contents[14'h0837] = 8'h68;
s_mem_contents[14'h0838] = 8'h08;
s_mem_contents[14'h0839] = 8'hc9;
s_mem_contents[14'h083a] = 8'hff;
s_mem_contents[14'h083b] = 8'hd0;
s_mem_contents[14'h083c] = 8'hfe;
s_mem_contents[14'h083d] = 8'h68;
s_mem_contents[14'h083e] = 8'h48;
s_mem_contents[14'h083f] = 8'hc9;
s_mem_contents[14'h0840] = 8'hb0;
s_mem_contents[14'h0841] = 8'hd0;
s_mem_contents[14'h0842] = 8'hfe;
s_mem_contents[14'h0843] = 8'h28;
s_mem_contents[14'h0844] = 8'ha9;
s_mem_contents[14'h0845] = 8'hff;
s_mem_contents[14'h0846] = 8'h48;
s_mem_contents[14'h0847] = 8'ha9;
s_mem_contents[14'h0848] = 8'hff;
s_mem_contents[14'h0849] = 8'h28;
s_mem_contents[14'h084a] = 8'h68;
s_mem_contents[14'h084b] = 8'h08;
s_mem_contents[14'h084c] = 8'hc9;
s_mem_contents[14'h084d] = 8'h00;
s_mem_contents[14'h084e] = 8'hd0;
s_mem_contents[14'h084f] = 8'hfe;
s_mem_contents[14'h0850] = 8'h68;
s_mem_contents[14'h0851] = 8'h48;
s_mem_contents[14'h0852] = 8'hc9;
s_mem_contents[14'h0853] = 8'h7f;
s_mem_contents[14'h0854] = 8'hd0;
s_mem_contents[14'h0855] = 8'hfe;
s_mem_contents[14'h0856] = 8'h28;
s_mem_contents[14'h0857] = 8'ha9;
s_mem_contents[14'h0858] = 8'h00;
s_mem_contents[14'h0859] = 8'h48;
s_mem_contents[14'h085a] = 8'ha9;
s_mem_contents[14'h085b] = 8'hfe;
s_mem_contents[14'h085c] = 8'h28;
s_mem_contents[14'h085d] = 8'h68;
s_mem_contents[14'h085e] = 8'h08;
s_mem_contents[14'h085f] = 8'hc9;
s_mem_contents[14'h0860] = 8'h01;
s_mem_contents[14'h0861] = 8'hd0;
s_mem_contents[14'h0862] = 8'hfe;
s_mem_contents[14'h0863] = 8'h68;
s_mem_contents[14'h0864] = 8'h48;
s_mem_contents[14'h0865] = 8'hc9;
s_mem_contents[14'h0866] = 8'h30;
s_mem_contents[14'h0867] = 8'hd0;
s_mem_contents[14'h0868] = 8'hfe;
s_mem_contents[14'h0869] = 8'h28;
s_mem_contents[14'h086a] = 8'he0;
s_mem_contents[14'h086b] = 8'h55;
s_mem_contents[14'h086c] = 8'hd0;
s_mem_contents[14'h086d] = 8'hfe;
s_mem_contents[14'h086e] = 8'hc0;
s_mem_contents[14'h086f] = 8'haa;
s_mem_contents[14'h0870] = 8'hd0;
s_mem_contents[14'h0871] = 8'hfe;
s_mem_contents[14'h0872] = 8'had;
s_mem_contents[14'h0873] = 8'h00;
s_mem_contents[14'h0874] = 8'h02;
s_mem_contents[14'h0875] = 8'hc9;
s_mem_contents[14'h0876] = 8'h05;
s_mem_contents[14'h0877] = 8'hd0;
s_mem_contents[14'h0878] = 8'hfe;
s_mem_contents[14'h0879] = 8'ha9;
s_mem_contents[14'h087a] = 8'h06;
s_mem_contents[14'h087b] = 8'h8d;
s_mem_contents[14'h087c] = 8'h00;
s_mem_contents[14'h087d] = 8'h02;
s_mem_contents[14'h087e] = 8'ha9;
s_mem_contents[14'h087f] = 8'h00;
s_mem_contents[14'h0880] = 8'h48;
s_mem_contents[14'h0881] = 8'ha9;
s_mem_contents[14'h0882] = 8'h3c;
s_mem_contents[14'h0883] = 8'h28;
s_mem_contents[14'h0884] = 8'h49;
s_mem_contents[14'h0885] = 8'hc3;
s_mem_contents[14'h0886] = 8'h08;
s_mem_contents[14'h0887] = 8'hc9;
s_mem_contents[14'h0888] = 8'hff;
s_mem_contents[14'h0889] = 8'hd0;
s_mem_contents[14'h088a] = 8'hfe;
s_mem_contents[14'h088b] = 8'h68;
s_mem_contents[14'h088c] = 8'h48;
s_mem_contents[14'h088d] = 8'hc9;
s_mem_contents[14'h088e] = 8'hb0;
s_mem_contents[14'h088f] = 8'hd0;
s_mem_contents[14'h0890] = 8'hfe;
s_mem_contents[14'h0891] = 8'h28;
s_mem_contents[14'h0892] = 8'ha9;
s_mem_contents[14'h0893] = 8'h00;
s_mem_contents[14'h0894] = 8'h48;
s_mem_contents[14'h0895] = 8'ha9;
s_mem_contents[14'h0896] = 8'hc3;
s_mem_contents[14'h0897] = 8'h28;
s_mem_contents[14'h0898] = 8'h49;
s_mem_contents[14'h0899] = 8'hc3;
s_mem_contents[14'h089a] = 8'h08;
s_mem_contents[14'h089b] = 8'hc9;
s_mem_contents[14'h089c] = 8'h00;
s_mem_contents[14'h089d] = 8'hd0;
s_mem_contents[14'h089e] = 8'hfe;
s_mem_contents[14'h089f] = 8'h68;
s_mem_contents[14'h08a0] = 8'h48;
s_mem_contents[14'h08a1] = 8'hc9;
s_mem_contents[14'h08a2] = 8'h32;
s_mem_contents[14'h08a3] = 8'hd0;
s_mem_contents[14'h08a4] = 8'hfe;
s_mem_contents[14'h08a5] = 8'h28;
s_mem_contents[14'h08a6] = 8'had;
s_mem_contents[14'h08a7] = 8'h00;
s_mem_contents[14'h08a8] = 8'h02;
s_mem_contents[14'h08a9] = 8'hc9;
s_mem_contents[14'h08aa] = 8'h06;
s_mem_contents[14'h08ab] = 8'hd0;
s_mem_contents[14'h08ac] = 8'hfe;
s_mem_contents[14'h08ad] = 8'ha9;
s_mem_contents[14'h08ae] = 8'h07;
s_mem_contents[14'h08af] = 8'h8d;
s_mem_contents[14'h08b0] = 8'h00;
s_mem_contents[14'h08b1] = 8'h02;
s_mem_contents[14'h08b2] = 8'ha2;
s_mem_contents[14'h08b3] = 8'h24;
s_mem_contents[14'h08b4] = 8'ha0;
s_mem_contents[14'h08b5] = 8'h42;
s_mem_contents[14'h08b6] = 8'ha9;
s_mem_contents[14'h08b7] = 8'h00;
s_mem_contents[14'h08b8] = 8'h48;
s_mem_contents[14'h08b9] = 8'ha9;
s_mem_contents[14'h08ba] = 8'h18;
s_mem_contents[14'h08bb] = 8'h28;
s_mem_contents[14'h08bc] = 8'hea;
s_mem_contents[14'h08bd] = 8'h08;
s_mem_contents[14'h08be] = 8'hc9;
s_mem_contents[14'h08bf] = 8'h18;
s_mem_contents[14'h08c0] = 8'hd0;
s_mem_contents[14'h08c1] = 8'hfe;
s_mem_contents[14'h08c2] = 8'h68;
s_mem_contents[14'h08c3] = 8'h48;
s_mem_contents[14'h08c4] = 8'hc9;
s_mem_contents[14'h08c5] = 8'h30;
s_mem_contents[14'h08c6] = 8'hd0;
s_mem_contents[14'h08c7] = 8'hfe;
s_mem_contents[14'h08c8] = 8'h28;
s_mem_contents[14'h08c9] = 8'he0;
s_mem_contents[14'h08ca] = 8'h24;
s_mem_contents[14'h08cb] = 8'hd0;
s_mem_contents[14'h08cc] = 8'hfe;
s_mem_contents[14'h08cd] = 8'hc0;
s_mem_contents[14'h08ce] = 8'h42;
s_mem_contents[14'h08cf] = 8'hd0;
s_mem_contents[14'h08d0] = 8'hfe;
s_mem_contents[14'h08d1] = 8'ha2;
s_mem_contents[14'h08d2] = 8'hdb;
s_mem_contents[14'h08d3] = 8'ha0;
s_mem_contents[14'h08d4] = 8'hbd;
s_mem_contents[14'h08d5] = 8'ha9;
s_mem_contents[14'h08d6] = 8'hff;
s_mem_contents[14'h08d7] = 8'h48;
s_mem_contents[14'h08d8] = 8'ha9;
s_mem_contents[14'h08d9] = 8'he7;
s_mem_contents[14'h08da] = 8'h28;
s_mem_contents[14'h08db] = 8'hea;
s_mem_contents[14'h08dc] = 8'h08;
s_mem_contents[14'h08dd] = 8'hc9;
s_mem_contents[14'h08de] = 8'he7;
s_mem_contents[14'h08df] = 8'hd0;
s_mem_contents[14'h08e0] = 8'hfe;
s_mem_contents[14'h08e1] = 8'h68;
s_mem_contents[14'h08e2] = 8'h48;
s_mem_contents[14'h08e3] = 8'hc9;
s_mem_contents[14'h08e4] = 8'hff;
s_mem_contents[14'h08e5] = 8'hd0;
s_mem_contents[14'h08e6] = 8'hfe;
s_mem_contents[14'h08e7] = 8'h28;
s_mem_contents[14'h08e8] = 8'he0;
s_mem_contents[14'h08e9] = 8'hdb;
s_mem_contents[14'h08ea] = 8'hd0;
s_mem_contents[14'h08eb] = 8'hfe;
s_mem_contents[14'h08ec] = 8'hc0;
s_mem_contents[14'h08ed] = 8'hbd;
s_mem_contents[14'h08ee] = 8'hd0;
s_mem_contents[14'h08ef] = 8'hfe;
s_mem_contents[14'h08f0] = 8'had;
s_mem_contents[14'h08f1] = 8'h00;
s_mem_contents[14'h08f2] = 8'h02;
s_mem_contents[14'h08f3] = 8'hc9;
s_mem_contents[14'h08f4] = 8'h07;
s_mem_contents[14'h08f5] = 8'hd0;
s_mem_contents[14'h08f6] = 8'hfe;
s_mem_contents[14'h08f7] = 8'ha9;
s_mem_contents[14'h08f8] = 8'h08;
s_mem_contents[14'h08f9] = 8'h8d;
s_mem_contents[14'h08fa] = 8'h00;
s_mem_contents[14'h08fb] = 8'h02;
s_mem_contents[14'h08fc] = 8'ha9;
s_mem_contents[14'h08fd] = 8'h00;
s_mem_contents[14'h08fe] = 8'h48;
s_mem_contents[14'h08ff] = 8'h28;
s_mem_contents[14'h0900] = 8'ha9;
s_mem_contents[14'h0901] = 8'h46;
s_mem_contents[14'h0902] = 8'ha2;
s_mem_contents[14'h0903] = 8'h41;
s_mem_contents[14'h0904] = 8'ha0;
s_mem_contents[14'h0905] = 8'h52;
s_mem_contents[14'h0906] = 8'h4c;
s_mem_contents[14'h0907] = 8'h74;
s_mem_contents[14'h0908] = 8'h34;
s_mem_contents[14'h0909] = 8'hea;
s_mem_contents[14'h090a] = 8'hea;
s_mem_contents[14'h090b] = 8'hd0;
s_mem_contents[14'h090c] = 8'hfe;
s_mem_contents[14'h090d] = 8'he8;
s_mem_contents[14'h090e] = 8'he8;
s_mem_contents[14'h090f] = 8'hf0;
s_mem_contents[14'h0910] = 8'hfe;
s_mem_contents[14'h0911] = 8'h10;
s_mem_contents[14'h0912] = 8'hfe;
s_mem_contents[14'h0913] = 8'h90;
s_mem_contents[14'h0914] = 8'hfe;
s_mem_contents[14'h0915] = 8'h50;
s_mem_contents[14'h0916] = 8'hfe;
s_mem_contents[14'h0917] = 8'hc9;
s_mem_contents[14'h0918] = 8'hec;
s_mem_contents[14'h0919] = 8'hd0;
s_mem_contents[14'h091a] = 8'hfe;
s_mem_contents[14'h091b] = 8'he0;
s_mem_contents[14'h091c] = 8'h42;
s_mem_contents[14'h091d] = 8'hd0;
s_mem_contents[14'h091e] = 8'hfe;
s_mem_contents[14'h091f] = 8'hc0;
s_mem_contents[14'h0920] = 8'h4f;
s_mem_contents[14'h0921] = 8'hd0;
s_mem_contents[14'h0922] = 8'hfe;
s_mem_contents[14'h0923] = 8'hca;
s_mem_contents[14'h0924] = 8'hc8;
s_mem_contents[14'h0925] = 8'hc8;
s_mem_contents[14'h0926] = 8'hc8;
s_mem_contents[14'h0927] = 8'h49;
s_mem_contents[14'h0928] = 8'haa;
s_mem_contents[14'h0929] = 8'h4c;
s_mem_contents[14'h092a] = 8'h32;
s_mem_contents[14'h092b] = 8'h09;
s_mem_contents[14'h092c] = 8'hea;
s_mem_contents[14'h092d] = 8'hea;
s_mem_contents[14'h092e] = 8'hd0;
s_mem_contents[14'h092f] = 8'hfe;
s_mem_contents[14'h0930] = 8'he8;
s_mem_contents[14'h0931] = 8'he8;
s_mem_contents[14'h0932] = 8'hf0;
s_mem_contents[14'h0933] = 8'hfe;
s_mem_contents[14'h0934] = 8'h30;
s_mem_contents[14'h0935] = 8'hfe;
s_mem_contents[14'h0936] = 8'h90;
s_mem_contents[14'h0937] = 8'hfe;
s_mem_contents[14'h0938] = 8'h50;
s_mem_contents[14'h0939] = 8'hfe;
s_mem_contents[14'h093a] = 8'hc9;
s_mem_contents[14'h093b] = 8'h46;
s_mem_contents[14'h093c] = 8'hd0;
s_mem_contents[14'h093d] = 8'hfe;
s_mem_contents[14'h093e] = 8'he0;
s_mem_contents[14'h093f] = 8'h41;
s_mem_contents[14'h0940] = 8'hd0;
s_mem_contents[14'h0941] = 8'hfe;
s_mem_contents[14'h0942] = 8'hc0;
s_mem_contents[14'h0943] = 8'h52;
s_mem_contents[14'h0944] = 8'hd0;
s_mem_contents[14'h0945] = 8'hfe;
s_mem_contents[14'h0946] = 8'had;
s_mem_contents[14'h0947] = 8'h00;
s_mem_contents[14'h0948] = 8'h02;
s_mem_contents[14'h0949] = 8'hc9;
s_mem_contents[14'h094a] = 8'h08;
s_mem_contents[14'h094b] = 8'hd0;
s_mem_contents[14'h094c] = 8'hfe;
s_mem_contents[14'h094d] = 8'ha9;
s_mem_contents[14'h094e] = 8'h09;
s_mem_contents[14'h094f] = 8'h8d;
s_mem_contents[14'h0950] = 8'h00;
s_mem_contents[14'h0951] = 8'h02;
s_mem_contents[14'h0952] = 8'ha9;
s_mem_contents[14'h0953] = 8'h00;
s_mem_contents[14'h0954] = 8'h48;
s_mem_contents[14'h0955] = 8'h28;
s_mem_contents[14'h0956] = 8'ha9;
s_mem_contents[14'h0957] = 8'h49;
s_mem_contents[14'h0958] = 8'ha2;
s_mem_contents[14'h0959] = 8'h4e;
s_mem_contents[14'h095a] = 8'ha0;
s_mem_contents[14'h095b] = 8'h44;
s_mem_contents[14'h095c] = 8'h6c;
s_mem_contents[14'h095d] = 8'ha2;
s_mem_contents[14'h095e] = 8'h34;
s_mem_contents[14'h095f] = 8'hea;
s_mem_contents[14'h0960] = 8'hd0;
s_mem_contents[14'h0961] = 8'hfe;
s_mem_contents[14'h0962] = 8'h88;
s_mem_contents[14'h0963] = 8'h88;
s_mem_contents[14'h0964] = 8'h08;
s_mem_contents[14'h0965] = 8'h88;
s_mem_contents[14'h0966] = 8'h88;
s_mem_contents[14'h0967] = 8'h88;
s_mem_contents[14'h0968] = 8'h28;
s_mem_contents[14'h0969] = 8'hf0;
s_mem_contents[14'h096a] = 8'hfe;
s_mem_contents[14'h096b] = 8'h10;
s_mem_contents[14'h096c] = 8'hfe;
s_mem_contents[14'h096d] = 8'h90;
s_mem_contents[14'h096e] = 8'hfe;
s_mem_contents[14'h096f] = 8'h50;
s_mem_contents[14'h0970] = 8'hfe;
s_mem_contents[14'h0971] = 8'hc9;
s_mem_contents[14'h0972] = 8'he3;
s_mem_contents[14'h0973] = 8'hd0;
s_mem_contents[14'h0974] = 8'hfe;
s_mem_contents[14'h0975] = 8'he0;
s_mem_contents[14'h0976] = 8'h4f;
s_mem_contents[14'h0977] = 8'hd0;
s_mem_contents[14'h0978] = 8'hfe;
s_mem_contents[14'h0979] = 8'hc0;
s_mem_contents[14'h097a] = 8'h3e;
s_mem_contents[14'h097b] = 8'hd0;
s_mem_contents[14'h097c] = 8'hfe;
s_mem_contents[14'h097d] = 8'hba;
s_mem_contents[14'h097e] = 8'he0;
s_mem_contents[14'h097f] = 8'hff;
s_mem_contents[14'h0980] = 8'hd0;
s_mem_contents[14'h0981] = 8'hfe;
s_mem_contents[14'h0982] = 8'had;
s_mem_contents[14'h0983] = 8'h00;
s_mem_contents[14'h0984] = 8'h02;
s_mem_contents[14'h0985] = 8'hc9;
s_mem_contents[14'h0986] = 8'h09;
s_mem_contents[14'h0987] = 8'hd0;
s_mem_contents[14'h0988] = 8'hfe;
s_mem_contents[14'h0989] = 8'ha9;
s_mem_contents[14'h098a] = 8'h0a;
s_mem_contents[14'h098b] = 8'h8d;
s_mem_contents[14'h098c] = 8'h00;
s_mem_contents[14'h098d] = 8'h02;
s_mem_contents[14'h098e] = 8'ha9;
s_mem_contents[14'h098f] = 8'h00;
s_mem_contents[14'h0990] = 8'h48;
s_mem_contents[14'h0991] = 8'h28;
s_mem_contents[14'h0992] = 8'ha9;
s_mem_contents[14'h0993] = 8'h4a;
s_mem_contents[14'h0994] = 8'ha2;
s_mem_contents[14'h0995] = 8'h53;
s_mem_contents[14'h0996] = 8'ha0;
s_mem_contents[14'h0997] = 8'h52;
s_mem_contents[14'h0998] = 8'h20;
s_mem_contents[14'h0999] = 8'he1;
s_mem_contents[14'h099a] = 8'h34;
s_mem_contents[14'h099b] = 8'h08;
s_mem_contents[14'h099c] = 8'h88;
s_mem_contents[14'h099d] = 8'h88;
s_mem_contents[14'h099e] = 8'h88;
s_mem_contents[14'h099f] = 8'h28;
s_mem_contents[14'h09a0] = 8'hf0;
s_mem_contents[14'h09a1] = 8'hfe;
s_mem_contents[14'h09a2] = 8'h10;
s_mem_contents[14'h09a3] = 8'hfe;
s_mem_contents[14'h09a4] = 8'h90;
s_mem_contents[14'h09a5] = 8'hfe;
s_mem_contents[14'h09a6] = 8'h50;
s_mem_contents[14'h09a7] = 8'hfe;
s_mem_contents[14'h09a8] = 8'hc9;
s_mem_contents[14'h09a9] = 8'he0;
s_mem_contents[14'h09aa] = 8'hd0;
s_mem_contents[14'h09ab] = 8'hfe;
s_mem_contents[14'h09ac] = 8'he0;
s_mem_contents[14'h09ad] = 8'h54;
s_mem_contents[14'h09ae] = 8'hd0;
s_mem_contents[14'h09af] = 8'hfe;
s_mem_contents[14'h09b0] = 8'hc0;
s_mem_contents[14'h09b1] = 8'h4c;
s_mem_contents[14'h09b2] = 8'hd0;
s_mem_contents[14'h09b3] = 8'hfe;
s_mem_contents[14'h09b4] = 8'hba;
s_mem_contents[14'h09b5] = 8'he0;
s_mem_contents[14'h09b6] = 8'hff;
s_mem_contents[14'h09b7] = 8'hd0;
s_mem_contents[14'h09b8] = 8'hfe;
s_mem_contents[14'h09b9] = 8'had;
s_mem_contents[14'h09ba] = 8'h00;
s_mem_contents[14'h09bb] = 8'h02;
s_mem_contents[14'h09bc] = 8'hc9;
s_mem_contents[14'h09bd] = 8'h0a;
s_mem_contents[14'h09be] = 8'hd0;
s_mem_contents[14'h09bf] = 8'hfe;
s_mem_contents[14'h09c0] = 8'ha9;
s_mem_contents[14'h09c1] = 8'h0b;
s_mem_contents[14'h09c2] = 8'h8d;
s_mem_contents[14'h09c3] = 8'h00;
s_mem_contents[14'h09c4] = 8'h02;
s_mem_contents[14'h09c5] = 8'had;
s_mem_contents[14'h09c6] = 8'h00;
s_mem_contents[14'h09c7] = 8'h02;
s_mem_contents[14'h09c8] = 8'hc9;
s_mem_contents[14'h09c9] = 8'h0b;
s_mem_contents[14'h09ca] = 8'hd0;
s_mem_contents[14'h09cb] = 8'hfe;
s_mem_contents[14'h09cc] = 8'ha9;
s_mem_contents[14'h09cd] = 8'h0c;
s_mem_contents[14'h09ce] = 8'h8d;
s_mem_contents[14'h09cf] = 8'h00;
s_mem_contents[14'h09d0] = 8'h02;
s_mem_contents[14'h09d1] = 8'ha9;
s_mem_contents[14'h09d2] = 8'hff;
s_mem_contents[14'h09d3] = 8'h48;
s_mem_contents[14'h09d4] = 8'h28;
s_mem_contents[14'h09d5] = 8'h18;
s_mem_contents[14'h09d6] = 8'h08;
s_mem_contents[14'h09d7] = 8'h68;
s_mem_contents[14'h09d8] = 8'h48;
s_mem_contents[14'h09d9] = 8'hc9;
s_mem_contents[14'h09da] = 8'hfe;
s_mem_contents[14'h09db] = 8'hd0;
s_mem_contents[14'h09dc] = 8'hfe;
s_mem_contents[14'h09dd] = 8'h28;
s_mem_contents[14'h09de] = 8'h38;
s_mem_contents[14'h09df] = 8'h08;
s_mem_contents[14'h09e0] = 8'h68;
s_mem_contents[14'h09e1] = 8'h48;
s_mem_contents[14'h09e2] = 8'hc9;
s_mem_contents[14'h09e3] = 8'hff;
s_mem_contents[14'h09e4] = 8'hd0;
s_mem_contents[14'h09e5] = 8'hfe;
s_mem_contents[14'h09e6] = 8'h28;
s_mem_contents[14'h09e7] = 8'h58;
s_mem_contents[14'h09e8] = 8'h08;
s_mem_contents[14'h09e9] = 8'h68;
s_mem_contents[14'h09ea] = 8'h48;
s_mem_contents[14'h09eb] = 8'hc9;
s_mem_contents[14'h09ec] = 8'hfb;
s_mem_contents[14'h09ed] = 8'hd0;
s_mem_contents[14'h09ee] = 8'hfe;
s_mem_contents[14'h09ef] = 8'h28;
s_mem_contents[14'h09f0] = 8'h78;
s_mem_contents[14'h09f1] = 8'h08;
s_mem_contents[14'h09f2] = 8'h68;
s_mem_contents[14'h09f3] = 8'h48;
s_mem_contents[14'h09f4] = 8'hc9;
s_mem_contents[14'h09f5] = 8'hff;
s_mem_contents[14'h09f6] = 8'hd0;
s_mem_contents[14'h09f7] = 8'hfe;
s_mem_contents[14'h09f8] = 8'h28;
s_mem_contents[14'h09f9] = 8'hd8;
s_mem_contents[14'h09fa] = 8'h08;
s_mem_contents[14'h09fb] = 8'h68;
s_mem_contents[14'h09fc] = 8'h48;
s_mem_contents[14'h09fd] = 8'hc9;
s_mem_contents[14'h09fe] = 8'hf7;
s_mem_contents[14'h09ff] = 8'hd0;
s_mem_contents[14'h0a00] = 8'hfe;
s_mem_contents[14'h0a01] = 8'h28;
s_mem_contents[14'h0a02] = 8'hf8;
s_mem_contents[14'h0a03] = 8'h08;
s_mem_contents[14'h0a04] = 8'h68;
s_mem_contents[14'h0a05] = 8'h48;
s_mem_contents[14'h0a06] = 8'hc9;
s_mem_contents[14'h0a07] = 8'hff;
s_mem_contents[14'h0a08] = 8'hd0;
s_mem_contents[14'h0a09] = 8'hfe;
s_mem_contents[14'h0a0a] = 8'h28;
s_mem_contents[14'h0a0b] = 8'hb8;
s_mem_contents[14'h0a0c] = 8'h08;
s_mem_contents[14'h0a0d] = 8'h68;
s_mem_contents[14'h0a0e] = 8'h48;
s_mem_contents[14'h0a0f] = 8'hc9;
s_mem_contents[14'h0a10] = 8'hbf;
s_mem_contents[14'h0a11] = 8'hd0;
s_mem_contents[14'h0a12] = 8'hfe;
s_mem_contents[14'h0a13] = 8'h28;
s_mem_contents[14'h0a14] = 8'ha9;
s_mem_contents[14'h0a15] = 8'h00;
s_mem_contents[14'h0a16] = 8'h48;
s_mem_contents[14'h0a17] = 8'h28;
s_mem_contents[14'h0a18] = 8'h08;
s_mem_contents[14'h0a19] = 8'h68;
s_mem_contents[14'h0a1a] = 8'h48;
s_mem_contents[14'h0a1b] = 8'hc9;
s_mem_contents[14'h0a1c] = 8'h30;
s_mem_contents[14'h0a1d] = 8'hd0;
s_mem_contents[14'h0a1e] = 8'hfe;
s_mem_contents[14'h0a1f] = 8'h28;
s_mem_contents[14'h0a20] = 8'h38;
s_mem_contents[14'h0a21] = 8'h08;
s_mem_contents[14'h0a22] = 8'h68;
s_mem_contents[14'h0a23] = 8'h48;
s_mem_contents[14'h0a24] = 8'hc9;
s_mem_contents[14'h0a25] = 8'h31;
s_mem_contents[14'h0a26] = 8'hd0;
s_mem_contents[14'h0a27] = 8'hfe;
s_mem_contents[14'h0a28] = 8'h28;
s_mem_contents[14'h0a29] = 8'h18;
s_mem_contents[14'h0a2a] = 8'h08;
s_mem_contents[14'h0a2b] = 8'h68;
s_mem_contents[14'h0a2c] = 8'h48;
s_mem_contents[14'h0a2d] = 8'hc9;
s_mem_contents[14'h0a2e] = 8'h30;
s_mem_contents[14'h0a2f] = 8'hd0;
s_mem_contents[14'h0a30] = 8'hfe;
s_mem_contents[14'h0a31] = 8'h28;
s_mem_contents[14'h0a32] = 8'h78;
s_mem_contents[14'h0a33] = 8'h08;
s_mem_contents[14'h0a34] = 8'h68;
s_mem_contents[14'h0a35] = 8'h48;
s_mem_contents[14'h0a36] = 8'hc9;
s_mem_contents[14'h0a37] = 8'h34;
s_mem_contents[14'h0a38] = 8'hd0;
s_mem_contents[14'h0a39] = 8'hfe;
s_mem_contents[14'h0a3a] = 8'h28;
s_mem_contents[14'h0a3b] = 8'h58;
s_mem_contents[14'h0a3c] = 8'h08;
s_mem_contents[14'h0a3d] = 8'h68;
s_mem_contents[14'h0a3e] = 8'h48;
s_mem_contents[14'h0a3f] = 8'hc9;
s_mem_contents[14'h0a40] = 8'h30;
s_mem_contents[14'h0a41] = 8'hd0;
s_mem_contents[14'h0a42] = 8'hfe;
s_mem_contents[14'h0a43] = 8'h28;
s_mem_contents[14'h0a44] = 8'hf8;
s_mem_contents[14'h0a45] = 8'h08;
s_mem_contents[14'h0a46] = 8'h68;
s_mem_contents[14'h0a47] = 8'h48;
s_mem_contents[14'h0a48] = 8'hc9;
s_mem_contents[14'h0a49] = 8'h38;
s_mem_contents[14'h0a4a] = 8'hd0;
s_mem_contents[14'h0a4b] = 8'hfe;
s_mem_contents[14'h0a4c] = 8'h28;
s_mem_contents[14'h0a4d] = 8'hd8;
s_mem_contents[14'h0a4e] = 8'h08;
s_mem_contents[14'h0a4f] = 8'h68;
s_mem_contents[14'h0a50] = 8'h48;
s_mem_contents[14'h0a51] = 8'hc9;
s_mem_contents[14'h0a52] = 8'h30;
s_mem_contents[14'h0a53] = 8'hd0;
s_mem_contents[14'h0a54] = 8'hfe;
s_mem_contents[14'h0a55] = 8'h28;
s_mem_contents[14'h0a56] = 8'ha9;
s_mem_contents[14'h0a57] = 8'h40;
s_mem_contents[14'h0a58] = 8'h48;
s_mem_contents[14'h0a59] = 8'h28;
s_mem_contents[14'h0a5a] = 8'h08;
s_mem_contents[14'h0a5b] = 8'h68;
s_mem_contents[14'h0a5c] = 8'h48;
s_mem_contents[14'h0a5d] = 8'hc9;
s_mem_contents[14'h0a5e] = 8'h70;
s_mem_contents[14'h0a5f] = 8'hd0;
s_mem_contents[14'h0a60] = 8'hfe;
s_mem_contents[14'h0a61] = 8'h28;
s_mem_contents[14'h0a62] = 8'hb8;
s_mem_contents[14'h0a63] = 8'h08;
s_mem_contents[14'h0a64] = 8'h68;
s_mem_contents[14'h0a65] = 8'h48;
s_mem_contents[14'h0a66] = 8'hc9;
s_mem_contents[14'h0a67] = 8'h30;
s_mem_contents[14'h0a68] = 8'hd0;
s_mem_contents[14'h0a69] = 8'hfe;
s_mem_contents[14'h0a6a] = 8'h28;
s_mem_contents[14'h0a6b] = 8'had;
s_mem_contents[14'h0a6c] = 8'h00;
s_mem_contents[14'h0a6d] = 8'h02;
s_mem_contents[14'h0a6e] = 8'hc9;
s_mem_contents[14'h0a6f] = 8'h0c;
s_mem_contents[14'h0a70] = 8'hd0;
s_mem_contents[14'h0a71] = 8'hfe;
s_mem_contents[14'h0a72] = 8'ha9;
s_mem_contents[14'h0a73] = 8'h0d;
s_mem_contents[14'h0a74] = 8'h8d;
s_mem_contents[14'h0a75] = 8'h00;
s_mem_contents[14'h0a76] = 8'h02;
s_mem_contents[14'h0a77] = 8'ha2;
s_mem_contents[14'h0a78] = 8'hfe;
s_mem_contents[14'h0a79] = 8'ha9;
s_mem_contents[14'h0a7a] = 8'hff;
s_mem_contents[14'h0a7b] = 8'h48;
s_mem_contents[14'h0a7c] = 8'h28;
s_mem_contents[14'h0a7d] = 8'he8;
s_mem_contents[14'h0a7e] = 8'h08;
s_mem_contents[14'h0a7f] = 8'he0;
s_mem_contents[14'h0a80] = 8'hff;
s_mem_contents[14'h0a81] = 8'hd0;
s_mem_contents[14'h0a82] = 8'hfe;
s_mem_contents[14'h0a83] = 8'h68;
s_mem_contents[14'h0a84] = 8'h48;
s_mem_contents[14'h0a85] = 8'hc9;
s_mem_contents[14'h0a86] = 8'hfd;
s_mem_contents[14'h0a87] = 8'hd0;
s_mem_contents[14'h0a88] = 8'hfe;
s_mem_contents[14'h0a89] = 8'h28;
s_mem_contents[14'h0a8a] = 8'he8;
s_mem_contents[14'h0a8b] = 8'h08;
s_mem_contents[14'h0a8c] = 8'he0;
s_mem_contents[14'h0a8d] = 8'h00;
s_mem_contents[14'h0a8e] = 8'hd0;
s_mem_contents[14'h0a8f] = 8'hfe;
s_mem_contents[14'h0a90] = 8'h68;
s_mem_contents[14'h0a91] = 8'h48;
s_mem_contents[14'h0a92] = 8'hc9;
s_mem_contents[14'h0a93] = 8'h7f;
s_mem_contents[14'h0a94] = 8'hd0;
s_mem_contents[14'h0a95] = 8'hfe;
s_mem_contents[14'h0a96] = 8'h28;
s_mem_contents[14'h0a97] = 8'he8;
s_mem_contents[14'h0a98] = 8'h08;
s_mem_contents[14'h0a99] = 8'he0;
s_mem_contents[14'h0a9a] = 8'h01;
s_mem_contents[14'h0a9b] = 8'hd0;
s_mem_contents[14'h0a9c] = 8'hfe;
s_mem_contents[14'h0a9d] = 8'h68;
s_mem_contents[14'h0a9e] = 8'h48;
s_mem_contents[14'h0a9f] = 8'hc9;
s_mem_contents[14'h0aa0] = 8'h7d;
s_mem_contents[14'h0aa1] = 8'hd0;
s_mem_contents[14'h0aa2] = 8'hfe;
s_mem_contents[14'h0aa3] = 8'h28;
s_mem_contents[14'h0aa4] = 8'hca;
s_mem_contents[14'h0aa5] = 8'h08;
s_mem_contents[14'h0aa6] = 8'he0;
s_mem_contents[14'h0aa7] = 8'h00;
s_mem_contents[14'h0aa8] = 8'hd0;
s_mem_contents[14'h0aa9] = 8'hfe;
s_mem_contents[14'h0aaa] = 8'h68;
s_mem_contents[14'h0aab] = 8'h48;
s_mem_contents[14'h0aac] = 8'hc9;
s_mem_contents[14'h0aad] = 8'h7f;
s_mem_contents[14'h0aae] = 8'hd0;
s_mem_contents[14'h0aaf] = 8'hfe;
s_mem_contents[14'h0ab0] = 8'h28;
s_mem_contents[14'h0ab1] = 8'hca;
s_mem_contents[14'h0ab2] = 8'h08;
s_mem_contents[14'h0ab3] = 8'he0;
s_mem_contents[14'h0ab4] = 8'hff;
s_mem_contents[14'h0ab5] = 8'hd0;
s_mem_contents[14'h0ab6] = 8'hfe;
s_mem_contents[14'h0ab7] = 8'h68;
s_mem_contents[14'h0ab8] = 8'h48;
s_mem_contents[14'h0ab9] = 8'hc9;
s_mem_contents[14'h0aba] = 8'hfd;
s_mem_contents[14'h0abb] = 8'hd0;
s_mem_contents[14'h0abc] = 8'hfe;
s_mem_contents[14'h0abd] = 8'h28;
s_mem_contents[14'h0abe] = 8'hca;
s_mem_contents[14'h0abf] = 8'ha9;
s_mem_contents[14'h0ac0] = 8'h00;
s_mem_contents[14'h0ac1] = 8'h48;
s_mem_contents[14'h0ac2] = 8'h28;
s_mem_contents[14'h0ac3] = 8'he8;
s_mem_contents[14'h0ac4] = 8'h08;
s_mem_contents[14'h0ac5] = 8'he0;
s_mem_contents[14'h0ac6] = 8'hff;
s_mem_contents[14'h0ac7] = 8'hd0;
s_mem_contents[14'h0ac8] = 8'hfe;
s_mem_contents[14'h0ac9] = 8'h68;
s_mem_contents[14'h0aca] = 8'h48;
s_mem_contents[14'h0acb] = 8'hc9;
s_mem_contents[14'h0acc] = 8'hb0;
s_mem_contents[14'h0acd] = 8'hd0;
s_mem_contents[14'h0ace] = 8'hfe;
s_mem_contents[14'h0acf] = 8'h28;
s_mem_contents[14'h0ad0] = 8'he8;
s_mem_contents[14'h0ad1] = 8'h08;
s_mem_contents[14'h0ad2] = 8'he0;
s_mem_contents[14'h0ad3] = 8'h00;
s_mem_contents[14'h0ad4] = 8'hd0;
s_mem_contents[14'h0ad5] = 8'hfe;
s_mem_contents[14'h0ad6] = 8'h68;
s_mem_contents[14'h0ad7] = 8'h48;
s_mem_contents[14'h0ad8] = 8'hc9;
s_mem_contents[14'h0ad9] = 8'h32;
s_mem_contents[14'h0ada] = 8'hd0;
s_mem_contents[14'h0adb] = 8'hfe;
s_mem_contents[14'h0adc] = 8'h28;
s_mem_contents[14'h0add] = 8'he8;
s_mem_contents[14'h0ade] = 8'h08;
s_mem_contents[14'h0adf] = 8'he0;
s_mem_contents[14'h0ae0] = 8'h01;
s_mem_contents[14'h0ae1] = 8'hd0;
s_mem_contents[14'h0ae2] = 8'hfe;
s_mem_contents[14'h0ae3] = 8'h68;
s_mem_contents[14'h0ae4] = 8'h48;
s_mem_contents[14'h0ae5] = 8'hc9;
s_mem_contents[14'h0ae6] = 8'h30;
s_mem_contents[14'h0ae7] = 8'hd0;
s_mem_contents[14'h0ae8] = 8'hfe;
s_mem_contents[14'h0ae9] = 8'h28;
s_mem_contents[14'h0aea] = 8'hca;
s_mem_contents[14'h0aeb] = 8'h08;
s_mem_contents[14'h0aec] = 8'he0;
s_mem_contents[14'h0aed] = 8'h00;
s_mem_contents[14'h0aee] = 8'hd0;
s_mem_contents[14'h0aef] = 8'hfe;
s_mem_contents[14'h0af0] = 8'h68;
s_mem_contents[14'h0af1] = 8'h48;
s_mem_contents[14'h0af2] = 8'hc9;
s_mem_contents[14'h0af3] = 8'h32;
s_mem_contents[14'h0af4] = 8'hd0;
s_mem_contents[14'h0af5] = 8'hfe;
s_mem_contents[14'h0af6] = 8'h28;
s_mem_contents[14'h0af7] = 8'hca;
s_mem_contents[14'h0af8] = 8'h08;
s_mem_contents[14'h0af9] = 8'he0;
s_mem_contents[14'h0afa] = 8'hff;
s_mem_contents[14'h0afb] = 8'hd0;
s_mem_contents[14'h0afc] = 8'hfe;
s_mem_contents[14'h0afd] = 8'h68;
s_mem_contents[14'h0afe] = 8'h48;
s_mem_contents[14'h0aff] = 8'hc9;
s_mem_contents[14'h0b00] = 8'hb0;
s_mem_contents[14'h0b01] = 8'hd0;
s_mem_contents[14'h0b02] = 8'hfe;
s_mem_contents[14'h0b03] = 8'h28;
s_mem_contents[14'h0b04] = 8'ha0;
s_mem_contents[14'h0b05] = 8'hfe;
s_mem_contents[14'h0b06] = 8'ha9;
s_mem_contents[14'h0b07] = 8'hff;
s_mem_contents[14'h0b08] = 8'h48;
s_mem_contents[14'h0b09] = 8'h28;
s_mem_contents[14'h0b0a] = 8'hc8;
s_mem_contents[14'h0b0b] = 8'h08;
s_mem_contents[14'h0b0c] = 8'hc0;
s_mem_contents[14'h0b0d] = 8'hff;
s_mem_contents[14'h0b0e] = 8'hd0;
s_mem_contents[14'h0b0f] = 8'hfe;
s_mem_contents[14'h0b10] = 8'h68;
s_mem_contents[14'h0b11] = 8'h48;
s_mem_contents[14'h0b12] = 8'hc9;
s_mem_contents[14'h0b13] = 8'hfd;
s_mem_contents[14'h0b14] = 8'hd0;
s_mem_contents[14'h0b15] = 8'hfe;
s_mem_contents[14'h0b16] = 8'h28;
s_mem_contents[14'h0b17] = 8'hc8;
s_mem_contents[14'h0b18] = 8'h08;
s_mem_contents[14'h0b19] = 8'hc0;
s_mem_contents[14'h0b1a] = 8'h00;
s_mem_contents[14'h0b1b] = 8'hd0;
s_mem_contents[14'h0b1c] = 8'hfe;
s_mem_contents[14'h0b1d] = 8'h68;
s_mem_contents[14'h0b1e] = 8'h48;
s_mem_contents[14'h0b1f] = 8'hc9;
s_mem_contents[14'h0b20] = 8'h7f;
s_mem_contents[14'h0b21] = 8'hd0;
s_mem_contents[14'h0b22] = 8'hfe;
s_mem_contents[14'h0b23] = 8'h28;
s_mem_contents[14'h0b24] = 8'hc8;
s_mem_contents[14'h0b25] = 8'h08;
s_mem_contents[14'h0b26] = 8'hc0;
s_mem_contents[14'h0b27] = 8'h01;
s_mem_contents[14'h0b28] = 8'hd0;
s_mem_contents[14'h0b29] = 8'hfe;
s_mem_contents[14'h0b2a] = 8'h68;
s_mem_contents[14'h0b2b] = 8'h48;
s_mem_contents[14'h0b2c] = 8'hc9;
s_mem_contents[14'h0b2d] = 8'h7d;
s_mem_contents[14'h0b2e] = 8'hd0;
s_mem_contents[14'h0b2f] = 8'hfe;
s_mem_contents[14'h0b30] = 8'h28;
s_mem_contents[14'h0b31] = 8'h88;
s_mem_contents[14'h0b32] = 8'h08;
s_mem_contents[14'h0b33] = 8'hc0;
s_mem_contents[14'h0b34] = 8'h00;
s_mem_contents[14'h0b35] = 8'hd0;
s_mem_contents[14'h0b36] = 8'hfe;
s_mem_contents[14'h0b37] = 8'h68;
s_mem_contents[14'h0b38] = 8'h48;
s_mem_contents[14'h0b39] = 8'hc9;
s_mem_contents[14'h0b3a] = 8'h7f;
s_mem_contents[14'h0b3b] = 8'hd0;
s_mem_contents[14'h0b3c] = 8'hfe;
s_mem_contents[14'h0b3d] = 8'h28;
s_mem_contents[14'h0b3e] = 8'h88;
s_mem_contents[14'h0b3f] = 8'h08;
s_mem_contents[14'h0b40] = 8'hc0;
s_mem_contents[14'h0b41] = 8'hff;
s_mem_contents[14'h0b42] = 8'hd0;
s_mem_contents[14'h0b43] = 8'hfe;
s_mem_contents[14'h0b44] = 8'h68;
s_mem_contents[14'h0b45] = 8'h48;
s_mem_contents[14'h0b46] = 8'hc9;
s_mem_contents[14'h0b47] = 8'hfd;
s_mem_contents[14'h0b48] = 8'hd0;
s_mem_contents[14'h0b49] = 8'hfe;
s_mem_contents[14'h0b4a] = 8'h28;
s_mem_contents[14'h0b4b] = 8'h88;
s_mem_contents[14'h0b4c] = 8'ha9;
s_mem_contents[14'h0b4d] = 8'h00;
s_mem_contents[14'h0b4e] = 8'h48;
s_mem_contents[14'h0b4f] = 8'h28;
s_mem_contents[14'h0b50] = 8'hc8;
s_mem_contents[14'h0b51] = 8'h08;
s_mem_contents[14'h0b52] = 8'hc0;
s_mem_contents[14'h0b53] = 8'hff;
s_mem_contents[14'h0b54] = 8'hd0;
s_mem_contents[14'h0b55] = 8'hfe;
s_mem_contents[14'h0b56] = 8'h68;
s_mem_contents[14'h0b57] = 8'h48;
s_mem_contents[14'h0b58] = 8'hc9;
s_mem_contents[14'h0b59] = 8'hb0;
s_mem_contents[14'h0b5a] = 8'hd0;
s_mem_contents[14'h0b5b] = 8'hfe;
s_mem_contents[14'h0b5c] = 8'h28;
s_mem_contents[14'h0b5d] = 8'hc8;
s_mem_contents[14'h0b5e] = 8'h08;
s_mem_contents[14'h0b5f] = 8'hc0;
s_mem_contents[14'h0b60] = 8'h00;
s_mem_contents[14'h0b61] = 8'hd0;
s_mem_contents[14'h0b62] = 8'hfe;
s_mem_contents[14'h0b63] = 8'h68;
s_mem_contents[14'h0b64] = 8'h48;
s_mem_contents[14'h0b65] = 8'hc9;
s_mem_contents[14'h0b66] = 8'h32;
s_mem_contents[14'h0b67] = 8'hd0;
s_mem_contents[14'h0b68] = 8'hfe;
s_mem_contents[14'h0b69] = 8'h28;
s_mem_contents[14'h0b6a] = 8'hc8;
s_mem_contents[14'h0b6b] = 8'h08;
s_mem_contents[14'h0b6c] = 8'hc0;
s_mem_contents[14'h0b6d] = 8'h01;
s_mem_contents[14'h0b6e] = 8'hd0;
s_mem_contents[14'h0b6f] = 8'hfe;
s_mem_contents[14'h0b70] = 8'h68;
s_mem_contents[14'h0b71] = 8'h48;
s_mem_contents[14'h0b72] = 8'hc9;
s_mem_contents[14'h0b73] = 8'h30;
s_mem_contents[14'h0b74] = 8'hd0;
s_mem_contents[14'h0b75] = 8'hfe;
s_mem_contents[14'h0b76] = 8'h28;
s_mem_contents[14'h0b77] = 8'h88;
s_mem_contents[14'h0b78] = 8'h08;
s_mem_contents[14'h0b79] = 8'hc0;
s_mem_contents[14'h0b7a] = 8'h00;
s_mem_contents[14'h0b7b] = 8'hd0;
s_mem_contents[14'h0b7c] = 8'hfe;
s_mem_contents[14'h0b7d] = 8'h68;
s_mem_contents[14'h0b7e] = 8'h48;
s_mem_contents[14'h0b7f] = 8'hc9;
s_mem_contents[14'h0b80] = 8'h32;
s_mem_contents[14'h0b81] = 8'hd0;
s_mem_contents[14'h0b82] = 8'hfe;
s_mem_contents[14'h0b83] = 8'h28;
s_mem_contents[14'h0b84] = 8'h88;
s_mem_contents[14'h0b85] = 8'h08;
s_mem_contents[14'h0b86] = 8'hc0;
s_mem_contents[14'h0b87] = 8'hff;
s_mem_contents[14'h0b88] = 8'hd0;
s_mem_contents[14'h0b89] = 8'hfe;
s_mem_contents[14'h0b8a] = 8'h68;
s_mem_contents[14'h0b8b] = 8'h48;
s_mem_contents[14'h0b8c] = 8'hc9;
s_mem_contents[14'h0b8d] = 8'hb0;
s_mem_contents[14'h0b8e] = 8'hd0;
s_mem_contents[14'h0b8f] = 8'hfe;
s_mem_contents[14'h0b90] = 8'h28;
s_mem_contents[14'h0b91] = 8'ha2;
s_mem_contents[14'h0b92] = 8'hff;
s_mem_contents[14'h0b93] = 8'ha9;
s_mem_contents[14'h0b94] = 8'hff;
s_mem_contents[14'h0b95] = 8'h48;
s_mem_contents[14'h0b96] = 8'h28;
s_mem_contents[14'h0b97] = 8'h8a;
s_mem_contents[14'h0b98] = 8'h08;
s_mem_contents[14'h0b99] = 8'hc9;
s_mem_contents[14'h0b9a] = 8'hff;
s_mem_contents[14'h0b9b] = 8'hd0;
s_mem_contents[14'h0b9c] = 8'hfe;
s_mem_contents[14'h0b9d] = 8'h68;
s_mem_contents[14'h0b9e] = 8'h48;
s_mem_contents[14'h0b9f] = 8'hc9;
s_mem_contents[14'h0ba0] = 8'hfd;
s_mem_contents[14'h0ba1] = 8'hd0;
s_mem_contents[14'h0ba2] = 8'hfe;
s_mem_contents[14'h0ba3] = 8'h28;
s_mem_contents[14'h0ba4] = 8'h08;
s_mem_contents[14'h0ba5] = 8'he8;
s_mem_contents[14'h0ba6] = 8'h28;
s_mem_contents[14'h0ba7] = 8'h8a;
s_mem_contents[14'h0ba8] = 8'h08;
s_mem_contents[14'h0ba9] = 8'hc9;
s_mem_contents[14'h0baa] = 8'h00;
s_mem_contents[14'h0bab] = 8'hd0;
s_mem_contents[14'h0bac] = 8'hfe;
s_mem_contents[14'h0bad] = 8'h68;
s_mem_contents[14'h0bae] = 8'h48;
s_mem_contents[14'h0baf] = 8'hc9;
s_mem_contents[14'h0bb0] = 8'h7f;
s_mem_contents[14'h0bb1] = 8'hd0;
s_mem_contents[14'h0bb2] = 8'hfe;
s_mem_contents[14'h0bb3] = 8'h28;
s_mem_contents[14'h0bb4] = 8'h08;
s_mem_contents[14'h0bb5] = 8'he8;
s_mem_contents[14'h0bb6] = 8'h28;
s_mem_contents[14'h0bb7] = 8'h8a;
s_mem_contents[14'h0bb8] = 8'h08;
s_mem_contents[14'h0bb9] = 8'hc9;
s_mem_contents[14'h0bba] = 8'h01;
s_mem_contents[14'h0bbb] = 8'hd0;
s_mem_contents[14'h0bbc] = 8'hfe;
s_mem_contents[14'h0bbd] = 8'h68;
s_mem_contents[14'h0bbe] = 8'h48;
s_mem_contents[14'h0bbf] = 8'hc9;
s_mem_contents[14'h0bc0] = 8'h7d;
s_mem_contents[14'h0bc1] = 8'hd0;
s_mem_contents[14'h0bc2] = 8'hfe;
s_mem_contents[14'h0bc3] = 8'h28;
s_mem_contents[14'h0bc4] = 8'ha9;
s_mem_contents[14'h0bc5] = 8'h00;
s_mem_contents[14'h0bc6] = 8'h48;
s_mem_contents[14'h0bc7] = 8'h28;
s_mem_contents[14'h0bc8] = 8'h8a;
s_mem_contents[14'h0bc9] = 8'h08;
s_mem_contents[14'h0bca] = 8'hc9;
s_mem_contents[14'h0bcb] = 8'h01;
s_mem_contents[14'h0bcc] = 8'hd0;
s_mem_contents[14'h0bcd] = 8'hfe;
s_mem_contents[14'h0bce] = 8'h68;
s_mem_contents[14'h0bcf] = 8'h48;
s_mem_contents[14'h0bd0] = 8'hc9;
s_mem_contents[14'h0bd1] = 8'h30;
s_mem_contents[14'h0bd2] = 8'hd0;
s_mem_contents[14'h0bd3] = 8'hfe;
s_mem_contents[14'h0bd4] = 8'h28;
s_mem_contents[14'h0bd5] = 8'h08;
s_mem_contents[14'h0bd6] = 8'hca;
s_mem_contents[14'h0bd7] = 8'h28;
s_mem_contents[14'h0bd8] = 8'h8a;
s_mem_contents[14'h0bd9] = 8'h08;
s_mem_contents[14'h0bda] = 8'hc9;
s_mem_contents[14'h0bdb] = 8'h00;
s_mem_contents[14'h0bdc] = 8'hd0;
s_mem_contents[14'h0bdd] = 8'hfe;
s_mem_contents[14'h0bde] = 8'h68;
s_mem_contents[14'h0bdf] = 8'h48;
s_mem_contents[14'h0be0] = 8'hc9;
s_mem_contents[14'h0be1] = 8'h32;
s_mem_contents[14'h0be2] = 8'hd0;
s_mem_contents[14'h0be3] = 8'hfe;
s_mem_contents[14'h0be4] = 8'h28;
s_mem_contents[14'h0be5] = 8'h08;
s_mem_contents[14'h0be6] = 8'hca;
s_mem_contents[14'h0be7] = 8'h28;
s_mem_contents[14'h0be8] = 8'h8a;
s_mem_contents[14'h0be9] = 8'h08;
s_mem_contents[14'h0bea] = 8'hc9;
s_mem_contents[14'h0beb] = 8'hff;
s_mem_contents[14'h0bec] = 8'hd0;
s_mem_contents[14'h0bed] = 8'hfe;
s_mem_contents[14'h0bee] = 8'h68;
s_mem_contents[14'h0bef] = 8'h48;
s_mem_contents[14'h0bf0] = 8'hc9;
s_mem_contents[14'h0bf1] = 8'hb0;
s_mem_contents[14'h0bf2] = 8'hd0;
s_mem_contents[14'h0bf3] = 8'hfe;
s_mem_contents[14'h0bf4] = 8'h28;
s_mem_contents[14'h0bf5] = 8'ha0;
s_mem_contents[14'h0bf6] = 8'hff;
s_mem_contents[14'h0bf7] = 8'ha9;
s_mem_contents[14'h0bf8] = 8'hff;
s_mem_contents[14'h0bf9] = 8'h48;
s_mem_contents[14'h0bfa] = 8'h28;
s_mem_contents[14'h0bfb] = 8'h98;
s_mem_contents[14'h0bfc] = 8'h08;
s_mem_contents[14'h0bfd] = 8'hc9;
s_mem_contents[14'h0bfe] = 8'hff;
s_mem_contents[14'h0bff] = 8'hd0;
s_mem_contents[14'h0c00] = 8'hfe;
s_mem_contents[14'h0c01] = 8'h68;
s_mem_contents[14'h0c02] = 8'h48;
s_mem_contents[14'h0c03] = 8'hc9;
s_mem_contents[14'h0c04] = 8'hfd;
s_mem_contents[14'h0c05] = 8'hd0;
s_mem_contents[14'h0c06] = 8'hfe;
s_mem_contents[14'h0c07] = 8'h28;
s_mem_contents[14'h0c08] = 8'h08;
s_mem_contents[14'h0c09] = 8'hc8;
s_mem_contents[14'h0c0a] = 8'h28;
s_mem_contents[14'h0c0b] = 8'h98;
s_mem_contents[14'h0c0c] = 8'h08;
s_mem_contents[14'h0c0d] = 8'hc9;
s_mem_contents[14'h0c0e] = 8'h00;
s_mem_contents[14'h0c0f] = 8'hd0;
s_mem_contents[14'h0c10] = 8'hfe;
s_mem_contents[14'h0c11] = 8'h68;
s_mem_contents[14'h0c12] = 8'h48;
s_mem_contents[14'h0c13] = 8'hc9;
s_mem_contents[14'h0c14] = 8'h7f;
s_mem_contents[14'h0c15] = 8'hd0;
s_mem_contents[14'h0c16] = 8'hfe;
s_mem_contents[14'h0c17] = 8'h28;
s_mem_contents[14'h0c18] = 8'h08;
s_mem_contents[14'h0c19] = 8'hc8;
s_mem_contents[14'h0c1a] = 8'h28;
s_mem_contents[14'h0c1b] = 8'h98;
s_mem_contents[14'h0c1c] = 8'h08;
s_mem_contents[14'h0c1d] = 8'hc9;
s_mem_contents[14'h0c1e] = 8'h01;
s_mem_contents[14'h0c1f] = 8'hd0;
s_mem_contents[14'h0c20] = 8'hfe;
s_mem_contents[14'h0c21] = 8'h68;
s_mem_contents[14'h0c22] = 8'h48;
s_mem_contents[14'h0c23] = 8'hc9;
s_mem_contents[14'h0c24] = 8'h7d;
s_mem_contents[14'h0c25] = 8'hd0;
s_mem_contents[14'h0c26] = 8'hfe;
s_mem_contents[14'h0c27] = 8'h28;
s_mem_contents[14'h0c28] = 8'ha9;
s_mem_contents[14'h0c29] = 8'h00;
s_mem_contents[14'h0c2a] = 8'h48;
s_mem_contents[14'h0c2b] = 8'h28;
s_mem_contents[14'h0c2c] = 8'h98;
s_mem_contents[14'h0c2d] = 8'h08;
s_mem_contents[14'h0c2e] = 8'hc9;
s_mem_contents[14'h0c2f] = 8'h01;
s_mem_contents[14'h0c30] = 8'hd0;
s_mem_contents[14'h0c31] = 8'hfe;
s_mem_contents[14'h0c32] = 8'h68;
s_mem_contents[14'h0c33] = 8'h48;
s_mem_contents[14'h0c34] = 8'hc9;
s_mem_contents[14'h0c35] = 8'h30;
s_mem_contents[14'h0c36] = 8'hd0;
s_mem_contents[14'h0c37] = 8'hfe;
s_mem_contents[14'h0c38] = 8'h28;
s_mem_contents[14'h0c39] = 8'h08;
s_mem_contents[14'h0c3a] = 8'h88;
s_mem_contents[14'h0c3b] = 8'h28;
s_mem_contents[14'h0c3c] = 8'h98;
s_mem_contents[14'h0c3d] = 8'h08;
s_mem_contents[14'h0c3e] = 8'hc9;
s_mem_contents[14'h0c3f] = 8'h00;
s_mem_contents[14'h0c40] = 8'hd0;
s_mem_contents[14'h0c41] = 8'hfe;
s_mem_contents[14'h0c42] = 8'h68;
s_mem_contents[14'h0c43] = 8'h48;
s_mem_contents[14'h0c44] = 8'hc9;
s_mem_contents[14'h0c45] = 8'h32;
s_mem_contents[14'h0c46] = 8'hd0;
s_mem_contents[14'h0c47] = 8'hfe;
s_mem_contents[14'h0c48] = 8'h28;
s_mem_contents[14'h0c49] = 8'h08;
s_mem_contents[14'h0c4a] = 8'h88;
s_mem_contents[14'h0c4b] = 8'h28;
s_mem_contents[14'h0c4c] = 8'h98;
s_mem_contents[14'h0c4d] = 8'h08;
s_mem_contents[14'h0c4e] = 8'hc9;
s_mem_contents[14'h0c4f] = 8'hff;
s_mem_contents[14'h0c50] = 8'hd0;
s_mem_contents[14'h0c51] = 8'hfe;
s_mem_contents[14'h0c52] = 8'h68;
s_mem_contents[14'h0c53] = 8'h48;
s_mem_contents[14'h0c54] = 8'hc9;
s_mem_contents[14'h0c55] = 8'hb0;
s_mem_contents[14'h0c56] = 8'hd0;
s_mem_contents[14'h0c57] = 8'hfe;
s_mem_contents[14'h0c58] = 8'h28;
s_mem_contents[14'h0c59] = 8'ha9;
s_mem_contents[14'h0c5a] = 8'hff;
s_mem_contents[14'h0c5b] = 8'h48;
s_mem_contents[14'h0c5c] = 8'ha2;
s_mem_contents[14'h0c5d] = 8'hff;
s_mem_contents[14'h0c5e] = 8'h8a;
s_mem_contents[14'h0c5f] = 8'h28;
s_mem_contents[14'h0c60] = 8'ha8;
s_mem_contents[14'h0c61] = 8'h08;
s_mem_contents[14'h0c62] = 8'hc0;
s_mem_contents[14'h0c63] = 8'hff;
s_mem_contents[14'h0c64] = 8'hd0;
s_mem_contents[14'h0c65] = 8'hfe;
s_mem_contents[14'h0c66] = 8'h68;
s_mem_contents[14'h0c67] = 8'h48;
s_mem_contents[14'h0c68] = 8'hc9;
s_mem_contents[14'h0c69] = 8'hfd;
s_mem_contents[14'h0c6a] = 8'hd0;
s_mem_contents[14'h0c6b] = 8'hfe;
s_mem_contents[14'h0c6c] = 8'h28;
s_mem_contents[14'h0c6d] = 8'h08;
s_mem_contents[14'h0c6e] = 8'he8;
s_mem_contents[14'h0c6f] = 8'h8a;
s_mem_contents[14'h0c70] = 8'h28;
s_mem_contents[14'h0c71] = 8'ha8;
s_mem_contents[14'h0c72] = 8'h08;
s_mem_contents[14'h0c73] = 8'hc0;
s_mem_contents[14'h0c74] = 8'h00;
s_mem_contents[14'h0c75] = 8'hd0;
s_mem_contents[14'h0c76] = 8'hfe;
s_mem_contents[14'h0c77] = 8'h68;
s_mem_contents[14'h0c78] = 8'h48;
s_mem_contents[14'h0c79] = 8'hc9;
s_mem_contents[14'h0c7a] = 8'h7f;
s_mem_contents[14'h0c7b] = 8'hd0;
s_mem_contents[14'h0c7c] = 8'hfe;
s_mem_contents[14'h0c7d] = 8'h28;
s_mem_contents[14'h0c7e] = 8'h08;
s_mem_contents[14'h0c7f] = 8'he8;
s_mem_contents[14'h0c80] = 8'h8a;
s_mem_contents[14'h0c81] = 8'h28;
s_mem_contents[14'h0c82] = 8'ha8;
s_mem_contents[14'h0c83] = 8'h08;
s_mem_contents[14'h0c84] = 8'hc0;
s_mem_contents[14'h0c85] = 8'h01;
s_mem_contents[14'h0c86] = 8'hd0;
s_mem_contents[14'h0c87] = 8'hfe;
s_mem_contents[14'h0c88] = 8'h68;
s_mem_contents[14'h0c89] = 8'h48;
s_mem_contents[14'h0c8a] = 8'hc9;
s_mem_contents[14'h0c8b] = 8'h7d;
s_mem_contents[14'h0c8c] = 8'hd0;
s_mem_contents[14'h0c8d] = 8'hfe;
s_mem_contents[14'h0c8e] = 8'h28;
s_mem_contents[14'h0c8f] = 8'ha9;
s_mem_contents[14'h0c90] = 8'h00;
s_mem_contents[14'h0c91] = 8'h48;
s_mem_contents[14'h0c92] = 8'ha9;
s_mem_contents[14'h0c93] = 8'h00;
s_mem_contents[14'h0c94] = 8'h8a;
s_mem_contents[14'h0c95] = 8'h28;
s_mem_contents[14'h0c96] = 8'ha8;
s_mem_contents[14'h0c97] = 8'h08;
s_mem_contents[14'h0c98] = 8'hc0;
s_mem_contents[14'h0c99] = 8'h01;
s_mem_contents[14'h0c9a] = 8'hd0;
s_mem_contents[14'h0c9b] = 8'hfe;
s_mem_contents[14'h0c9c] = 8'h68;
s_mem_contents[14'h0c9d] = 8'h48;
s_mem_contents[14'h0c9e] = 8'hc9;
s_mem_contents[14'h0c9f] = 8'h30;
s_mem_contents[14'h0ca0] = 8'hd0;
s_mem_contents[14'h0ca1] = 8'hfe;
s_mem_contents[14'h0ca2] = 8'h28;
s_mem_contents[14'h0ca3] = 8'h08;
s_mem_contents[14'h0ca4] = 8'hca;
s_mem_contents[14'h0ca5] = 8'h8a;
s_mem_contents[14'h0ca6] = 8'h28;
s_mem_contents[14'h0ca7] = 8'ha8;
s_mem_contents[14'h0ca8] = 8'h08;
s_mem_contents[14'h0ca9] = 8'hc0;
s_mem_contents[14'h0caa] = 8'h00;
s_mem_contents[14'h0cab] = 8'hd0;
s_mem_contents[14'h0cac] = 8'hfe;
s_mem_contents[14'h0cad] = 8'h68;
s_mem_contents[14'h0cae] = 8'h48;
s_mem_contents[14'h0caf] = 8'hc9;
s_mem_contents[14'h0cb0] = 8'h32;
s_mem_contents[14'h0cb1] = 8'hd0;
s_mem_contents[14'h0cb2] = 8'hfe;
s_mem_contents[14'h0cb3] = 8'h28;
s_mem_contents[14'h0cb4] = 8'h08;
s_mem_contents[14'h0cb5] = 8'hca;
s_mem_contents[14'h0cb6] = 8'h8a;
s_mem_contents[14'h0cb7] = 8'h28;
s_mem_contents[14'h0cb8] = 8'ha8;
s_mem_contents[14'h0cb9] = 8'h08;
s_mem_contents[14'h0cba] = 8'hc0;
s_mem_contents[14'h0cbb] = 8'hff;
s_mem_contents[14'h0cbc] = 8'hd0;
s_mem_contents[14'h0cbd] = 8'hfe;
s_mem_contents[14'h0cbe] = 8'h68;
s_mem_contents[14'h0cbf] = 8'h48;
s_mem_contents[14'h0cc0] = 8'hc9;
s_mem_contents[14'h0cc1] = 8'hb0;
s_mem_contents[14'h0cc2] = 8'hd0;
s_mem_contents[14'h0cc3] = 8'hfe;
s_mem_contents[14'h0cc4] = 8'h28;
s_mem_contents[14'h0cc5] = 8'ha9;
s_mem_contents[14'h0cc6] = 8'hff;
s_mem_contents[14'h0cc7] = 8'h48;
s_mem_contents[14'h0cc8] = 8'ha0;
s_mem_contents[14'h0cc9] = 8'hff;
s_mem_contents[14'h0cca] = 8'h98;
s_mem_contents[14'h0ccb] = 8'h28;
s_mem_contents[14'h0ccc] = 8'haa;
s_mem_contents[14'h0ccd] = 8'h08;
s_mem_contents[14'h0cce] = 8'he0;
s_mem_contents[14'h0ccf] = 8'hff;
s_mem_contents[14'h0cd0] = 8'hd0;
s_mem_contents[14'h0cd1] = 8'hfe;
s_mem_contents[14'h0cd2] = 8'h68;
s_mem_contents[14'h0cd3] = 8'h48;
s_mem_contents[14'h0cd4] = 8'hc9;
s_mem_contents[14'h0cd5] = 8'hfd;
s_mem_contents[14'h0cd6] = 8'hd0;
s_mem_contents[14'h0cd7] = 8'hfe;
s_mem_contents[14'h0cd8] = 8'h28;
s_mem_contents[14'h0cd9] = 8'h08;
s_mem_contents[14'h0cda] = 8'hc8;
s_mem_contents[14'h0cdb] = 8'h98;
s_mem_contents[14'h0cdc] = 8'h28;
s_mem_contents[14'h0cdd] = 8'haa;
s_mem_contents[14'h0cde] = 8'h08;
s_mem_contents[14'h0cdf] = 8'he0;
s_mem_contents[14'h0ce0] = 8'h00;
s_mem_contents[14'h0ce1] = 8'hd0;
s_mem_contents[14'h0ce2] = 8'hfe;
s_mem_contents[14'h0ce3] = 8'h68;
s_mem_contents[14'h0ce4] = 8'h48;
s_mem_contents[14'h0ce5] = 8'hc9;
s_mem_contents[14'h0ce6] = 8'h7f;
s_mem_contents[14'h0ce7] = 8'hd0;
s_mem_contents[14'h0ce8] = 8'hfe;
s_mem_contents[14'h0ce9] = 8'h28;
s_mem_contents[14'h0cea] = 8'h08;
s_mem_contents[14'h0ceb] = 8'hc8;
s_mem_contents[14'h0cec] = 8'h98;
s_mem_contents[14'h0ced] = 8'h28;
s_mem_contents[14'h0cee] = 8'haa;
s_mem_contents[14'h0cef] = 8'h08;
s_mem_contents[14'h0cf0] = 8'he0;
s_mem_contents[14'h0cf1] = 8'h01;
s_mem_contents[14'h0cf2] = 8'hd0;
s_mem_contents[14'h0cf3] = 8'hfe;
s_mem_contents[14'h0cf4] = 8'h68;
s_mem_contents[14'h0cf5] = 8'h48;
s_mem_contents[14'h0cf6] = 8'hc9;
s_mem_contents[14'h0cf7] = 8'h7d;
s_mem_contents[14'h0cf8] = 8'hd0;
s_mem_contents[14'h0cf9] = 8'hfe;
s_mem_contents[14'h0cfa] = 8'h28;
s_mem_contents[14'h0cfb] = 8'ha9;
s_mem_contents[14'h0cfc] = 8'h00;
s_mem_contents[14'h0cfd] = 8'h48;
s_mem_contents[14'h0cfe] = 8'ha9;
s_mem_contents[14'h0cff] = 8'h00;
s_mem_contents[14'h0d00] = 8'h98;
s_mem_contents[14'h0d01] = 8'h28;
s_mem_contents[14'h0d02] = 8'haa;
s_mem_contents[14'h0d03] = 8'h08;
s_mem_contents[14'h0d04] = 8'he0;
s_mem_contents[14'h0d05] = 8'h01;
s_mem_contents[14'h0d06] = 8'hd0;
s_mem_contents[14'h0d07] = 8'hfe;
s_mem_contents[14'h0d08] = 8'h68;
s_mem_contents[14'h0d09] = 8'h48;
s_mem_contents[14'h0d0a] = 8'hc9;
s_mem_contents[14'h0d0b] = 8'h30;
s_mem_contents[14'h0d0c] = 8'hd0;
s_mem_contents[14'h0d0d] = 8'hfe;
s_mem_contents[14'h0d0e] = 8'h28;
s_mem_contents[14'h0d0f] = 8'h08;
s_mem_contents[14'h0d10] = 8'h88;
s_mem_contents[14'h0d11] = 8'h98;
s_mem_contents[14'h0d12] = 8'h28;
s_mem_contents[14'h0d13] = 8'haa;
s_mem_contents[14'h0d14] = 8'h08;
s_mem_contents[14'h0d15] = 8'he0;
s_mem_contents[14'h0d16] = 8'h00;
s_mem_contents[14'h0d17] = 8'hd0;
s_mem_contents[14'h0d18] = 8'hfe;
s_mem_contents[14'h0d19] = 8'h68;
s_mem_contents[14'h0d1a] = 8'h48;
s_mem_contents[14'h0d1b] = 8'hc9;
s_mem_contents[14'h0d1c] = 8'h32;
s_mem_contents[14'h0d1d] = 8'hd0;
s_mem_contents[14'h0d1e] = 8'hfe;
s_mem_contents[14'h0d1f] = 8'h28;
s_mem_contents[14'h0d20] = 8'h08;
s_mem_contents[14'h0d21] = 8'h88;
s_mem_contents[14'h0d22] = 8'h98;
s_mem_contents[14'h0d23] = 8'h28;
s_mem_contents[14'h0d24] = 8'haa;
s_mem_contents[14'h0d25] = 8'h08;
s_mem_contents[14'h0d26] = 8'he0;
s_mem_contents[14'h0d27] = 8'hff;
s_mem_contents[14'h0d28] = 8'hd0;
s_mem_contents[14'h0d29] = 8'hfe;
s_mem_contents[14'h0d2a] = 8'h68;
s_mem_contents[14'h0d2b] = 8'h48;
s_mem_contents[14'h0d2c] = 8'hc9;
s_mem_contents[14'h0d2d] = 8'hb0;
s_mem_contents[14'h0d2e] = 8'hd0;
s_mem_contents[14'h0d2f] = 8'hfe;
s_mem_contents[14'h0d30] = 8'h28;
s_mem_contents[14'h0d31] = 8'had;
s_mem_contents[14'h0d32] = 8'h00;
s_mem_contents[14'h0d33] = 8'h02;
s_mem_contents[14'h0d34] = 8'hc9;
s_mem_contents[14'h0d35] = 8'h0d;
s_mem_contents[14'h0d36] = 8'hd0;
s_mem_contents[14'h0d37] = 8'hfe;
s_mem_contents[14'h0d38] = 8'ha9;
s_mem_contents[14'h0d39] = 8'h0e;
s_mem_contents[14'h0d3a] = 8'h8d;
s_mem_contents[14'h0d3b] = 8'h00;
s_mem_contents[14'h0d3c] = 8'h02;
s_mem_contents[14'h0d3d] = 8'ha2;
s_mem_contents[14'h0d3e] = 8'h01;
s_mem_contents[14'h0d3f] = 8'ha9;
s_mem_contents[14'h0d40] = 8'hff;
s_mem_contents[14'h0d41] = 8'h48;
s_mem_contents[14'h0d42] = 8'h28;
s_mem_contents[14'h0d43] = 8'h9a;
s_mem_contents[14'h0d44] = 8'h08;
s_mem_contents[14'h0d45] = 8'had;
s_mem_contents[14'h0d46] = 8'h01;
s_mem_contents[14'h0d47] = 8'h01;
s_mem_contents[14'h0d48] = 8'hc9;
s_mem_contents[14'h0d49] = 8'hff;
s_mem_contents[14'h0d4a] = 8'hd0;
s_mem_contents[14'h0d4b] = 8'hfe;
s_mem_contents[14'h0d4c] = 8'ha9;
s_mem_contents[14'h0d4d] = 8'h00;
s_mem_contents[14'h0d4e] = 8'h48;
s_mem_contents[14'h0d4f] = 8'h28;
s_mem_contents[14'h0d50] = 8'h9a;
s_mem_contents[14'h0d51] = 8'h08;
s_mem_contents[14'h0d52] = 8'had;
s_mem_contents[14'h0d53] = 8'h01;
s_mem_contents[14'h0d54] = 8'h01;
s_mem_contents[14'h0d55] = 8'hc9;
s_mem_contents[14'h0d56] = 8'h30;
s_mem_contents[14'h0d57] = 8'hd0;
s_mem_contents[14'h0d58] = 8'hfe;
s_mem_contents[14'h0d59] = 8'hca;
s_mem_contents[14'h0d5a] = 8'ha9;
s_mem_contents[14'h0d5b] = 8'hff;
s_mem_contents[14'h0d5c] = 8'h48;
s_mem_contents[14'h0d5d] = 8'h28;
s_mem_contents[14'h0d5e] = 8'h9a;
s_mem_contents[14'h0d5f] = 8'h08;
s_mem_contents[14'h0d60] = 8'had;
s_mem_contents[14'h0d61] = 8'h00;
s_mem_contents[14'h0d62] = 8'h01;
s_mem_contents[14'h0d63] = 8'hc9;
s_mem_contents[14'h0d64] = 8'hff;
s_mem_contents[14'h0d65] = 8'hd0;
s_mem_contents[14'h0d66] = 8'hfe;
s_mem_contents[14'h0d67] = 8'ha9;
s_mem_contents[14'h0d68] = 8'h00;
s_mem_contents[14'h0d69] = 8'h48;
s_mem_contents[14'h0d6a] = 8'h28;
s_mem_contents[14'h0d6b] = 8'h9a;
s_mem_contents[14'h0d6c] = 8'h08;
s_mem_contents[14'h0d6d] = 8'had;
s_mem_contents[14'h0d6e] = 8'h00;
s_mem_contents[14'h0d6f] = 8'h01;
s_mem_contents[14'h0d70] = 8'hc9;
s_mem_contents[14'h0d71] = 8'h30;
s_mem_contents[14'h0d72] = 8'hd0;
s_mem_contents[14'h0d73] = 8'hfe;
s_mem_contents[14'h0d74] = 8'hca;
s_mem_contents[14'h0d75] = 8'ha9;
s_mem_contents[14'h0d76] = 8'hff;
s_mem_contents[14'h0d77] = 8'h48;
s_mem_contents[14'h0d78] = 8'h28;
s_mem_contents[14'h0d79] = 8'h9a;
s_mem_contents[14'h0d7a] = 8'h08;
s_mem_contents[14'h0d7b] = 8'had;
s_mem_contents[14'h0d7c] = 8'hff;
s_mem_contents[14'h0d7d] = 8'h01;
s_mem_contents[14'h0d7e] = 8'hc9;
s_mem_contents[14'h0d7f] = 8'hff;
s_mem_contents[14'h0d80] = 8'hd0;
s_mem_contents[14'h0d81] = 8'hfe;
s_mem_contents[14'h0d82] = 8'ha9;
s_mem_contents[14'h0d83] = 8'h00;
s_mem_contents[14'h0d84] = 8'h48;
s_mem_contents[14'h0d85] = 8'h28;
s_mem_contents[14'h0d86] = 8'h9a;
s_mem_contents[14'h0d87] = 8'h08;
s_mem_contents[14'h0d88] = 8'had;
s_mem_contents[14'h0d89] = 8'hff;
s_mem_contents[14'h0d8a] = 8'h01;
s_mem_contents[14'h0d8b] = 8'hc9;
s_mem_contents[14'h0d8c] = 8'h30;
s_mem_contents[14'h0d8d] = 8'ha2;
s_mem_contents[14'h0d8e] = 8'h01;
s_mem_contents[14'h0d8f] = 8'h9a;
s_mem_contents[14'h0d90] = 8'ha9;
s_mem_contents[14'h0d91] = 8'hff;
s_mem_contents[14'h0d92] = 8'h48;
s_mem_contents[14'h0d93] = 8'h28;
s_mem_contents[14'h0d94] = 8'hba;
s_mem_contents[14'h0d95] = 8'h08;
s_mem_contents[14'h0d96] = 8'he0;
s_mem_contents[14'h0d97] = 8'h01;
s_mem_contents[14'h0d98] = 8'hd0;
s_mem_contents[14'h0d99] = 8'hfe;
s_mem_contents[14'h0d9a] = 8'had;
s_mem_contents[14'h0d9b] = 8'h01;
s_mem_contents[14'h0d9c] = 8'h01;
s_mem_contents[14'h0d9d] = 8'hc9;
s_mem_contents[14'h0d9e] = 8'h7d;
s_mem_contents[14'h0d9f] = 8'hd0;
s_mem_contents[14'h0da0] = 8'hfe;
s_mem_contents[14'h0da1] = 8'ha9;
s_mem_contents[14'h0da2] = 8'hff;
s_mem_contents[14'h0da3] = 8'h48;
s_mem_contents[14'h0da4] = 8'h28;
s_mem_contents[14'h0da5] = 8'hba;
s_mem_contents[14'h0da6] = 8'h08;
s_mem_contents[14'h0da7] = 8'he0;
s_mem_contents[14'h0da8] = 8'h00;
s_mem_contents[14'h0da9] = 8'hd0;
s_mem_contents[14'h0daa] = 8'hfe;
s_mem_contents[14'h0dab] = 8'had;
s_mem_contents[14'h0dac] = 8'h00;
s_mem_contents[14'h0dad] = 8'h01;
s_mem_contents[14'h0dae] = 8'hc9;
s_mem_contents[14'h0daf] = 8'h7f;
s_mem_contents[14'h0db0] = 8'hd0;
s_mem_contents[14'h0db1] = 8'hfe;
s_mem_contents[14'h0db2] = 8'ha9;
s_mem_contents[14'h0db3] = 8'hff;
s_mem_contents[14'h0db4] = 8'h48;
s_mem_contents[14'h0db5] = 8'h28;
s_mem_contents[14'h0db6] = 8'hba;
s_mem_contents[14'h0db7] = 8'h08;
s_mem_contents[14'h0db8] = 8'he0;
s_mem_contents[14'h0db9] = 8'hff;
s_mem_contents[14'h0dba] = 8'hd0;
s_mem_contents[14'h0dbb] = 8'hfe;
s_mem_contents[14'h0dbc] = 8'had;
s_mem_contents[14'h0dbd] = 8'hff;
s_mem_contents[14'h0dbe] = 8'h01;
s_mem_contents[14'h0dbf] = 8'hc9;
s_mem_contents[14'h0dc0] = 8'hfd;
s_mem_contents[14'h0dc1] = 8'hd0;
s_mem_contents[14'h0dc2] = 8'hfe;
s_mem_contents[14'h0dc3] = 8'ha2;
s_mem_contents[14'h0dc4] = 8'h01;
s_mem_contents[14'h0dc5] = 8'h9a;
s_mem_contents[14'h0dc6] = 8'ha9;
s_mem_contents[14'h0dc7] = 8'h00;
s_mem_contents[14'h0dc8] = 8'h48;
s_mem_contents[14'h0dc9] = 8'h28;
s_mem_contents[14'h0dca] = 8'hba;
s_mem_contents[14'h0dcb] = 8'h08;
s_mem_contents[14'h0dcc] = 8'he0;
s_mem_contents[14'h0dcd] = 8'h01;
s_mem_contents[14'h0dce] = 8'hd0;
s_mem_contents[14'h0dcf] = 8'hfe;
s_mem_contents[14'h0dd0] = 8'had;
s_mem_contents[14'h0dd1] = 8'h01;
s_mem_contents[14'h0dd2] = 8'h01;
s_mem_contents[14'h0dd3] = 8'hc9;
s_mem_contents[14'h0dd4] = 8'h30;
s_mem_contents[14'h0dd5] = 8'hd0;
s_mem_contents[14'h0dd6] = 8'hfe;
s_mem_contents[14'h0dd7] = 8'ha9;
s_mem_contents[14'h0dd8] = 8'h00;
s_mem_contents[14'h0dd9] = 8'h48;
s_mem_contents[14'h0dda] = 8'h28;
s_mem_contents[14'h0ddb] = 8'hba;
s_mem_contents[14'h0ddc] = 8'h08;
s_mem_contents[14'h0ddd] = 8'he0;
s_mem_contents[14'h0dde] = 8'h00;
s_mem_contents[14'h0ddf] = 8'hd0;
s_mem_contents[14'h0de0] = 8'hfe;
s_mem_contents[14'h0de1] = 8'had;
s_mem_contents[14'h0de2] = 8'h00;
s_mem_contents[14'h0de3] = 8'h01;
s_mem_contents[14'h0de4] = 8'hc9;
s_mem_contents[14'h0de5] = 8'h32;
s_mem_contents[14'h0de6] = 8'hd0;
s_mem_contents[14'h0de7] = 8'hfe;
s_mem_contents[14'h0de8] = 8'ha9;
s_mem_contents[14'h0de9] = 8'h00;
s_mem_contents[14'h0dea] = 8'h48;
s_mem_contents[14'h0deb] = 8'h28;
s_mem_contents[14'h0dec] = 8'hba;
s_mem_contents[14'h0ded] = 8'h08;
s_mem_contents[14'h0dee] = 8'he0;
s_mem_contents[14'h0def] = 8'hff;
s_mem_contents[14'h0df0] = 8'hd0;
s_mem_contents[14'h0df1] = 8'hfe;
s_mem_contents[14'h0df2] = 8'had;
s_mem_contents[14'h0df3] = 8'hff;
s_mem_contents[14'h0df4] = 8'h01;
s_mem_contents[14'h0df5] = 8'hc9;
s_mem_contents[14'h0df6] = 8'hb0;
s_mem_contents[14'h0df7] = 8'hd0;
s_mem_contents[14'h0df8] = 8'hfe;
s_mem_contents[14'h0df9] = 8'h68;
s_mem_contents[14'h0dfa] = 8'had;
s_mem_contents[14'h0dfb] = 8'h00;
s_mem_contents[14'h0dfc] = 8'h02;
s_mem_contents[14'h0dfd] = 8'hc9;
s_mem_contents[14'h0dfe] = 8'h0e;
s_mem_contents[14'h0dff] = 8'hd0;
s_mem_contents[14'h0e00] = 8'hfe;
s_mem_contents[14'h0e01] = 8'ha9;
s_mem_contents[14'h0e02] = 8'h0f;
s_mem_contents[14'h0e03] = 8'h8d;
s_mem_contents[14'h0e04] = 8'h00;
s_mem_contents[14'h0e05] = 8'h02;
s_mem_contents[14'h0e06] = 8'ha0;
s_mem_contents[14'h0e07] = 8'h03;
s_mem_contents[14'h0e08] = 8'ha9;
s_mem_contents[14'h0e09] = 8'h00;
s_mem_contents[14'h0e0a] = 8'h48;
s_mem_contents[14'h0e0b] = 8'h28;
s_mem_contents[14'h0e0c] = 8'hb6;
s_mem_contents[14'h0e0d] = 8'h09;
s_mem_contents[14'h0e0e] = 8'h08;
s_mem_contents[14'h0e0f] = 8'h8a;
s_mem_contents[14'h0e10] = 8'h49;
s_mem_contents[14'h0e11] = 8'hc3;
s_mem_contents[14'h0e12] = 8'h28;
s_mem_contents[14'h0e13] = 8'h99;
s_mem_contents[14'h0e14] = 8'h03;
s_mem_contents[14'h0e15] = 8'h02;
s_mem_contents[14'h0e16] = 8'h08;
s_mem_contents[14'h0e17] = 8'h49;
s_mem_contents[14'h0e18] = 8'hc3;
s_mem_contents[14'h0e19] = 8'hd9;
s_mem_contents[14'h0e1a] = 8'h17;
s_mem_contents[14'h0e1b] = 8'h02;
s_mem_contents[14'h0e1c] = 8'hd0;
s_mem_contents[14'h0e1d] = 8'hfe;
s_mem_contents[14'h0e1e] = 8'h68;
s_mem_contents[14'h0e1f] = 8'h49;
s_mem_contents[14'h0e20] = 8'h30;
s_mem_contents[14'h0e21] = 8'hd9;
s_mem_contents[14'h0e22] = 8'h1c;
s_mem_contents[14'h0e23] = 8'h02;
s_mem_contents[14'h0e24] = 8'hd0;
s_mem_contents[14'h0e25] = 8'hfe;
s_mem_contents[14'h0e26] = 8'h88;
s_mem_contents[14'h0e27] = 8'h10;
s_mem_contents[14'h0e28] = 8'hdf;
s_mem_contents[14'h0e29] = 8'ha0;
s_mem_contents[14'h0e2a] = 8'h03;
s_mem_contents[14'h0e2b] = 8'ha9;
s_mem_contents[14'h0e2c] = 8'hff;
s_mem_contents[14'h0e2d] = 8'h48;
s_mem_contents[14'h0e2e] = 8'h28;
s_mem_contents[14'h0e2f] = 8'hb6;
s_mem_contents[14'h0e30] = 8'h09;
s_mem_contents[14'h0e31] = 8'h08;
s_mem_contents[14'h0e32] = 8'h8a;
s_mem_contents[14'h0e33] = 8'h49;
s_mem_contents[14'h0e34] = 8'hc3;
s_mem_contents[14'h0e35] = 8'h28;
s_mem_contents[14'h0e36] = 8'h99;
s_mem_contents[14'h0e37] = 8'h03;
s_mem_contents[14'h0e38] = 8'h02;
s_mem_contents[14'h0e39] = 8'h08;
s_mem_contents[14'h0e3a] = 8'h49;
s_mem_contents[14'h0e3b] = 8'hc3;
s_mem_contents[14'h0e3c] = 8'hd9;
s_mem_contents[14'h0e3d] = 8'h17;
s_mem_contents[14'h0e3e] = 8'h02;
s_mem_contents[14'h0e3f] = 8'hd0;
s_mem_contents[14'h0e40] = 8'hfe;
s_mem_contents[14'h0e41] = 8'h68;
s_mem_contents[14'h0e42] = 8'h49;
s_mem_contents[14'h0e43] = 8'h7d;
s_mem_contents[14'h0e44] = 8'hd9;
s_mem_contents[14'h0e45] = 8'h1c;
s_mem_contents[14'h0e46] = 8'h02;
s_mem_contents[14'h0e47] = 8'hd0;
s_mem_contents[14'h0e48] = 8'hfe;
s_mem_contents[14'h0e49] = 8'h88;
s_mem_contents[14'h0e4a] = 8'h10;
s_mem_contents[14'h0e4b] = 8'hdf;
s_mem_contents[14'h0e4c] = 8'ha0;
s_mem_contents[14'h0e4d] = 8'h03;
s_mem_contents[14'h0e4e] = 8'ha9;
s_mem_contents[14'h0e4f] = 8'h00;
s_mem_contents[14'h0e50] = 8'h48;
s_mem_contents[14'h0e51] = 8'h28;
s_mem_contents[14'h0e52] = 8'hbe;
s_mem_contents[14'h0e53] = 8'h17;
s_mem_contents[14'h0e54] = 8'h02;
s_mem_contents[14'h0e55] = 8'h08;
s_mem_contents[14'h0e56] = 8'h8a;
s_mem_contents[14'h0e57] = 8'h49;
s_mem_contents[14'h0e58] = 8'hc3;
s_mem_contents[14'h0e59] = 8'haa;
s_mem_contents[14'h0e5a] = 8'h28;
s_mem_contents[14'h0e5b] = 8'h96;
s_mem_contents[14'h0e5c] = 8'h02;
s_mem_contents[14'h0e5d] = 8'h08;
s_mem_contents[14'h0e5e] = 8'h49;
s_mem_contents[14'h0e5f] = 8'hc3;
s_mem_contents[14'h0e60] = 8'hd9;
s_mem_contents[14'h0e61] = 8'h09;
s_mem_contents[14'h0e62] = 8'h00;
s_mem_contents[14'h0e63] = 8'hd0;
s_mem_contents[14'h0e64] = 8'hfe;
s_mem_contents[14'h0e65] = 8'h68;
s_mem_contents[14'h0e66] = 8'h49;
s_mem_contents[14'h0e67] = 8'h30;
s_mem_contents[14'h0e68] = 8'hd9;
s_mem_contents[14'h0e69] = 8'h1c;
s_mem_contents[14'h0e6a] = 8'h02;
s_mem_contents[14'h0e6b] = 8'hd0;
s_mem_contents[14'h0e6c] = 8'hfe;
s_mem_contents[14'h0e6d] = 8'h88;
s_mem_contents[14'h0e6e] = 8'h10;
s_mem_contents[14'h0e6f] = 8'hde;
s_mem_contents[14'h0e70] = 8'ha0;
s_mem_contents[14'h0e71] = 8'h03;
s_mem_contents[14'h0e72] = 8'ha9;
s_mem_contents[14'h0e73] = 8'hff;
s_mem_contents[14'h0e74] = 8'h48;
s_mem_contents[14'h0e75] = 8'h28;
s_mem_contents[14'h0e76] = 8'hbe;
s_mem_contents[14'h0e77] = 8'h17;
s_mem_contents[14'h0e78] = 8'h02;
s_mem_contents[14'h0e79] = 8'h08;
s_mem_contents[14'h0e7a] = 8'h8a;
s_mem_contents[14'h0e7b] = 8'h49;
s_mem_contents[14'h0e7c] = 8'hc3;
s_mem_contents[14'h0e7d] = 8'haa;
s_mem_contents[14'h0e7e] = 8'h28;
s_mem_contents[14'h0e7f] = 8'h96;
s_mem_contents[14'h0e80] = 8'h02;
s_mem_contents[14'h0e81] = 8'h08;
s_mem_contents[14'h0e82] = 8'h49;
s_mem_contents[14'h0e83] = 8'hc3;
s_mem_contents[14'h0e84] = 8'hd9;
s_mem_contents[14'h0e85] = 8'h09;
s_mem_contents[14'h0e86] = 8'h00;
s_mem_contents[14'h0e87] = 8'hd0;
s_mem_contents[14'h0e88] = 8'hfe;
s_mem_contents[14'h0e89] = 8'h68;
s_mem_contents[14'h0e8a] = 8'h49;
s_mem_contents[14'h0e8b] = 8'h7d;
s_mem_contents[14'h0e8c] = 8'hd9;
s_mem_contents[14'h0e8d] = 8'h1c;
s_mem_contents[14'h0e8e] = 8'h02;
s_mem_contents[14'h0e8f] = 8'hd0;
s_mem_contents[14'h0e90] = 8'hfe;
s_mem_contents[14'h0e91] = 8'h88;
s_mem_contents[14'h0e92] = 8'h10;
s_mem_contents[14'h0e93] = 8'hde;
s_mem_contents[14'h0e94] = 8'ha0;
s_mem_contents[14'h0e95] = 8'h03;
s_mem_contents[14'h0e96] = 8'ha2;
s_mem_contents[14'h0e97] = 8'h00;
s_mem_contents[14'h0e98] = 8'hb9;
s_mem_contents[14'h0e99] = 8'h02;
s_mem_contents[14'h0e9a] = 8'h00;
s_mem_contents[14'h0e9b] = 8'h49;
s_mem_contents[14'h0e9c] = 8'hc3;
s_mem_contents[14'h0e9d] = 8'hd9;
s_mem_contents[14'h0e9e] = 8'h09;
s_mem_contents[14'h0e9f] = 8'h00;
s_mem_contents[14'h0ea0] = 8'hd0;
s_mem_contents[14'h0ea1] = 8'hfe;
s_mem_contents[14'h0ea2] = 8'h96;
s_mem_contents[14'h0ea3] = 8'h02;
s_mem_contents[14'h0ea4] = 8'hb9;
s_mem_contents[14'h0ea5] = 8'h03;
s_mem_contents[14'h0ea6] = 8'h02;
s_mem_contents[14'h0ea7] = 8'h49;
s_mem_contents[14'h0ea8] = 8'hc3;
s_mem_contents[14'h0ea9] = 8'hd9;
s_mem_contents[14'h0eaa] = 8'h17;
s_mem_contents[14'h0eab] = 8'h02;
s_mem_contents[14'h0eac] = 8'hd0;
s_mem_contents[14'h0ead] = 8'hfe;
s_mem_contents[14'h0eae] = 8'h8a;
s_mem_contents[14'h0eaf] = 8'h99;
s_mem_contents[14'h0eb0] = 8'h03;
s_mem_contents[14'h0eb1] = 8'h02;
s_mem_contents[14'h0eb2] = 8'h88;
s_mem_contents[14'h0eb3] = 8'h10;
s_mem_contents[14'h0eb4] = 8'he3;
s_mem_contents[14'h0eb5] = 8'had;
s_mem_contents[14'h0eb6] = 8'h00;
s_mem_contents[14'h0eb7] = 8'h02;
s_mem_contents[14'h0eb8] = 8'hc9;
s_mem_contents[14'h0eb9] = 8'h0f;
s_mem_contents[14'h0eba] = 8'hd0;
s_mem_contents[14'h0ebb] = 8'hfe;
s_mem_contents[14'h0ebc] = 8'ha9;
s_mem_contents[14'h0ebd] = 8'h10;
s_mem_contents[14'h0ebe] = 8'h8d;
s_mem_contents[14'h0ebf] = 8'h00;
s_mem_contents[14'h0ec0] = 8'h02;
s_mem_contents[14'h0ec1] = 8'ha0;
s_mem_contents[14'h0ec2] = 8'hfd;
s_mem_contents[14'h0ec3] = 8'hb6;
s_mem_contents[14'h0ec4] = 8'h0f;
s_mem_contents[14'h0ec5] = 8'h8a;
s_mem_contents[14'h0ec6] = 8'h99;
s_mem_contents[14'h0ec7] = 8'h09;
s_mem_contents[14'h0ec8] = 8'h01;
s_mem_contents[14'h0ec9] = 8'h88;
s_mem_contents[14'h0eca] = 8'hc0;
s_mem_contents[14'h0ecb] = 8'hfa;
s_mem_contents[14'h0ecc] = 8'hb0;
s_mem_contents[14'h0ecd] = 8'hf5;
s_mem_contents[14'h0ece] = 8'ha0;
s_mem_contents[14'h0ecf] = 8'hfd;
s_mem_contents[14'h0ed0] = 8'hbe;
s_mem_contents[14'h0ed1] = 8'h1d;
s_mem_contents[14'h0ed2] = 8'h01;
s_mem_contents[14'h0ed3] = 8'h96;
s_mem_contents[14'h0ed4] = 8'h08;
s_mem_contents[14'h0ed5] = 8'h88;
s_mem_contents[14'h0ed6] = 8'hc0;
s_mem_contents[14'h0ed7] = 8'hfa;
s_mem_contents[14'h0ed8] = 8'hb0;
s_mem_contents[14'h0ed9] = 8'hf6;
s_mem_contents[14'h0eda] = 8'ha0;
s_mem_contents[14'h0edb] = 8'h03;
s_mem_contents[14'h0edc] = 8'ha2;
s_mem_contents[14'h0edd] = 8'h00;
s_mem_contents[14'h0ede] = 8'hb9;
s_mem_contents[14'h0edf] = 8'h02;
s_mem_contents[14'h0ee0] = 8'h00;
s_mem_contents[14'h0ee1] = 8'hd9;
s_mem_contents[14'h0ee2] = 8'h09;
s_mem_contents[14'h0ee3] = 8'h00;
s_mem_contents[14'h0ee4] = 8'hd0;
s_mem_contents[14'h0ee5] = 8'hfe;
s_mem_contents[14'h0ee6] = 8'h96;
s_mem_contents[14'h0ee7] = 8'h02;
s_mem_contents[14'h0ee8] = 8'hb9;
s_mem_contents[14'h0ee9] = 8'h03;
s_mem_contents[14'h0eea] = 8'h02;
s_mem_contents[14'h0eeb] = 8'hd9;
s_mem_contents[14'h0eec] = 8'h17;
s_mem_contents[14'h0eed] = 8'h02;
s_mem_contents[14'h0eee] = 8'hd0;
s_mem_contents[14'h0eef] = 8'hfe;
s_mem_contents[14'h0ef0] = 8'h8a;
s_mem_contents[14'h0ef1] = 8'h99;
s_mem_contents[14'h0ef2] = 8'h03;
s_mem_contents[14'h0ef3] = 8'h02;
s_mem_contents[14'h0ef4] = 8'h88;
s_mem_contents[14'h0ef5] = 8'h10;
s_mem_contents[14'h0ef6] = 8'he7;
s_mem_contents[14'h0ef7] = 8'had;
s_mem_contents[14'h0ef8] = 8'h00;
s_mem_contents[14'h0ef9] = 8'h02;
s_mem_contents[14'h0efa] = 8'hc9;
s_mem_contents[14'h0efb] = 8'h10;
s_mem_contents[14'h0efc] = 8'hd0;
s_mem_contents[14'h0efd] = 8'hfe;
s_mem_contents[14'h0efe] = 8'ha9;
s_mem_contents[14'h0eff] = 8'h11;
s_mem_contents[14'h0f00] = 8'h8d;
s_mem_contents[14'h0f01] = 8'h00;
s_mem_contents[14'h0f02] = 8'h02;
s_mem_contents[14'h0f03] = 8'ha2;
s_mem_contents[14'h0f04] = 8'h03;
s_mem_contents[14'h0f05] = 8'ha9;
s_mem_contents[14'h0f06] = 8'h00;
s_mem_contents[14'h0f07] = 8'h48;
s_mem_contents[14'h0f08] = 8'h28;
s_mem_contents[14'h0f09] = 8'hb4;
s_mem_contents[14'h0f0a] = 8'h09;
s_mem_contents[14'h0f0b] = 8'h08;
s_mem_contents[14'h0f0c] = 8'h98;
s_mem_contents[14'h0f0d] = 8'h49;
s_mem_contents[14'h0f0e] = 8'hc3;
s_mem_contents[14'h0f0f] = 8'h28;
s_mem_contents[14'h0f10] = 8'h9d;
s_mem_contents[14'h0f11] = 8'h03;
s_mem_contents[14'h0f12] = 8'h02;
s_mem_contents[14'h0f13] = 8'h08;
s_mem_contents[14'h0f14] = 8'h49;
s_mem_contents[14'h0f15] = 8'hc3;
s_mem_contents[14'h0f16] = 8'hdd;
s_mem_contents[14'h0f17] = 8'h17;
s_mem_contents[14'h0f18] = 8'h02;
s_mem_contents[14'h0f19] = 8'hd0;
s_mem_contents[14'h0f1a] = 8'hfe;
s_mem_contents[14'h0f1b] = 8'h68;
s_mem_contents[14'h0f1c] = 8'h49;
s_mem_contents[14'h0f1d] = 8'h30;
s_mem_contents[14'h0f1e] = 8'hdd;
s_mem_contents[14'h0f1f] = 8'h1c;
s_mem_contents[14'h0f20] = 8'h02;
s_mem_contents[14'h0f21] = 8'hd0;
s_mem_contents[14'h0f22] = 8'hfe;
s_mem_contents[14'h0f23] = 8'hca;
s_mem_contents[14'h0f24] = 8'h10;
s_mem_contents[14'h0f25] = 8'hdf;
s_mem_contents[14'h0f26] = 8'ha2;
s_mem_contents[14'h0f27] = 8'h03;
s_mem_contents[14'h0f28] = 8'ha9;
s_mem_contents[14'h0f29] = 8'hff;
s_mem_contents[14'h0f2a] = 8'h48;
s_mem_contents[14'h0f2b] = 8'h28;
s_mem_contents[14'h0f2c] = 8'hb4;
s_mem_contents[14'h0f2d] = 8'h09;
s_mem_contents[14'h0f2e] = 8'h08;
s_mem_contents[14'h0f2f] = 8'h98;
s_mem_contents[14'h0f30] = 8'h49;
s_mem_contents[14'h0f31] = 8'hc3;
s_mem_contents[14'h0f32] = 8'h28;
s_mem_contents[14'h0f33] = 8'h9d;
s_mem_contents[14'h0f34] = 8'h03;
s_mem_contents[14'h0f35] = 8'h02;
s_mem_contents[14'h0f36] = 8'h08;
s_mem_contents[14'h0f37] = 8'h49;
s_mem_contents[14'h0f38] = 8'hc3;
s_mem_contents[14'h0f39] = 8'hdd;
s_mem_contents[14'h0f3a] = 8'h17;
s_mem_contents[14'h0f3b] = 8'h02;
s_mem_contents[14'h0f3c] = 8'hd0;
s_mem_contents[14'h0f3d] = 8'hfe;
s_mem_contents[14'h0f3e] = 8'h68;
s_mem_contents[14'h0f3f] = 8'h49;
s_mem_contents[14'h0f40] = 8'h7d;
s_mem_contents[14'h0f41] = 8'hdd;
s_mem_contents[14'h0f42] = 8'h1c;
s_mem_contents[14'h0f43] = 8'h02;
s_mem_contents[14'h0f44] = 8'hd0;
s_mem_contents[14'h0f45] = 8'hfe;
s_mem_contents[14'h0f46] = 8'hca;
s_mem_contents[14'h0f47] = 8'h10;
s_mem_contents[14'h0f48] = 8'hdf;
s_mem_contents[14'h0f49] = 8'ha2;
s_mem_contents[14'h0f4a] = 8'h03;
s_mem_contents[14'h0f4b] = 8'ha9;
s_mem_contents[14'h0f4c] = 8'h00;
s_mem_contents[14'h0f4d] = 8'h48;
s_mem_contents[14'h0f4e] = 8'h28;
s_mem_contents[14'h0f4f] = 8'hbc;
s_mem_contents[14'h0f50] = 8'h17;
s_mem_contents[14'h0f51] = 8'h02;
s_mem_contents[14'h0f52] = 8'h08;
s_mem_contents[14'h0f53] = 8'h98;
s_mem_contents[14'h0f54] = 8'h49;
s_mem_contents[14'h0f55] = 8'hc3;
s_mem_contents[14'h0f56] = 8'ha8;
s_mem_contents[14'h0f57] = 8'h28;
s_mem_contents[14'h0f58] = 8'h94;
s_mem_contents[14'h0f59] = 8'h02;
s_mem_contents[14'h0f5a] = 8'h08;
s_mem_contents[14'h0f5b] = 8'h49;
s_mem_contents[14'h0f5c] = 8'hc3;
s_mem_contents[14'h0f5d] = 8'hd5;
s_mem_contents[14'h0f5e] = 8'h09;
s_mem_contents[14'h0f5f] = 8'hd0;
s_mem_contents[14'h0f60] = 8'hfe;
s_mem_contents[14'h0f61] = 8'h68;
s_mem_contents[14'h0f62] = 8'h49;
s_mem_contents[14'h0f63] = 8'h30;
s_mem_contents[14'h0f64] = 8'hdd;
s_mem_contents[14'h0f65] = 8'h1c;
s_mem_contents[14'h0f66] = 8'h02;
s_mem_contents[14'h0f67] = 8'hd0;
s_mem_contents[14'h0f68] = 8'hfe;
s_mem_contents[14'h0f69] = 8'hca;
s_mem_contents[14'h0f6a] = 8'h10;
s_mem_contents[14'h0f6b] = 8'hdf;
s_mem_contents[14'h0f6c] = 8'ha2;
s_mem_contents[14'h0f6d] = 8'h03;
s_mem_contents[14'h0f6e] = 8'ha9;
s_mem_contents[14'h0f6f] = 8'hff;
s_mem_contents[14'h0f70] = 8'h48;
s_mem_contents[14'h0f71] = 8'h28;
s_mem_contents[14'h0f72] = 8'hbc;
s_mem_contents[14'h0f73] = 8'h17;
s_mem_contents[14'h0f74] = 8'h02;
s_mem_contents[14'h0f75] = 8'h08;
s_mem_contents[14'h0f76] = 8'h98;
s_mem_contents[14'h0f77] = 8'h49;
s_mem_contents[14'h0f78] = 8'hc3;
s_mem_contents[14'h0f79] = 8'ha8;
s_mem_contents[14'h0f7a] = 8'h28;
s_mem_contents[14'h0f7b] = 8'h94;
s_mem_contents[14'h0f7c] = 8'h02;
s_mem_contents[14'h0f7d] = 8'h08;
s_mem_contents[14'h0f7e] = 8'h49;
s_mem_contents[14'h0f7f] = 8'hc3;
s_mem_contents[14'h0f80] = 8'hd5;
s_mem_contents[14'h0f81] = 8'h09;
s_mem_contents[14'h0f82] = 8'hd0;
s_mem_contents[14'h0f83] = 8'hfe;
s_mem_contents[14'h0f84] = 8'h68;
s_mem_contents[14'h0f85] = 8'h49;
s_mem_contents[14'h0f86] = 8'h7d;
s_mem_contents[14'h0f87] = 8'hdd;
s_mem_contents[14'h0f88] = 8'h1c;
s_mem_contents[14'h0f89] = 8'h02;
s_mem_contents[14'h0f8a] = 8'hd0;
s_mem_contents[14'h0f8b] = 8'hfe;
s_mem_contents[14'h0f8c] = 8'hca;
s_mem_contents[14'h0f8d] = 8'h10;
s_mem_contents[14'h0f8e] = 8'hdf;
s_mem_contents[14'h0f8f] = 8'ha2;
s_mem_contents[14'h0f90] = 8'h03;
s_mem_contents[14'h0f91] = 8'ha0;
s_mem_contents[14'h0f92] = 8'h00;
s_mem_contents[14'h0f93] = 8'hb5;
s_mem_contents[14'h0f94] = 8'h02;
s_mem_contents[14'h0f95] = 8'h49;
s_mem_contents[14'h0f96] = 8'hc3;
s_mem_contents[14'h0f97] = 8'hd5;
s_mem_contents[14'h0f98] = 8'h09;
s_mem_contents[14'h0f99] = 8'hd0;
s_mem_contents[14'h0f9a] = 8'hfe;
s_mem_contents[14'h0f9b] = 8'h94;
s_mem_contents[14'h0f9c] = 8'h02;
s_mem_contents[14'h0f9d] = 8'hbd;
s_mem_contents[14'h0f9e] = 8'h03;
s_mem_contents[14'h0f9f] = 8'h02;
s_mem_contents[14'h0fa0] = 8'h49;
s_mem_contents[14'h0fa1] = 8'hc3;
s_mem_contents[14'h0fa2] = 8'hdd;
s_mem_contents[14'h0fa3] = 8'h17;
s_mem_contents[14'h0fa4] = 8'h02;
s_mem_contents[14'h0fa5] = 8'hd0;
s_mem_contents[14'h0fa6] = 8'hfe;
s_mem_contents[14'h0fa7] = 8'h8a;
s_mem_contents[14'h0fa8] = 8'h9d;
s_mem_contents[14'h0fa9] = 8'h03;
s_mem_contents[14'h0faa] = 8'h02;
s_mem_contents[14'h0fab] = 8'hca;
s_mem_contents[14'h0fac] = 8'h10;
s_mem_contents[14'h0fad] = 8'he5;
s_mem_contents[14'h0fae] = 8'had;
s_mem_contents[14'h0faf] = 8'h00;
s_mem_contents[14'h0fb0] = 8'h02;
s_mem_contents[14'h0fb1] = 8'hc9;
s_mem_contents[14'h0fb2] = 8'h11;
s_mem_contents[14'h0fb3] = 8'hd0;
s_mem_contents[14'h0fb4] = 8'hfe;
s_mem_contents[14'h0fb5] = 8'ha9;
s_mem_contents[14'h0fb6] = 8'h12;
s_mem_contents[14'h0fb7] = 8'h8d;
s_mem_contents[14'h0fb8] = 8'h00;
s_mem_contents[14'h0fb9] = 8'h02;
s_mem_contents[14'h0fba] = 8'ha2;
s_mem_contents[14'h0fbb] = 8'hfd;
s_mem_contents[14'h0fbc] = 8'hb4;
s_mem_contents[14'h0fbd] = 8'h0f;
s_mem_contents[14'h0fbe] = 8'h98;
s_mem_contents[14'h0fbf] = 8'h9d;
s_mem_contents[14'h0fc0] = 8'h09;
s_mem_contents[14'h0fc1] = 8'h01;
s_mem_contents[14'h0fc2] = 8'hca;
s_mem_contents[14'h0fc3] = 8'he0;
s_mem_contents[14'h0fc4] = 8'hfa;
s_mem_contents[14'h0fc5] = 8'hb0;
s_mem_contents[14'h0fc6] = 8'hf5;
s_mem_contents[14'h0fc7] = 8'ha2;
s_mem_contents[14'h0fc8] = 8'hfd;
s_mem_contents[14'h0fc9] = 8'hbc;
s_mem_contents[14'h0fca] = 8'h1d;
s_mem_contents[14'h0fcb] = 8'h01;
s_mem_contents[14'h0fcc] = 8'h94;
s_mem_contents[14'h0fcd] = 8'h08;
s_mem_contents[14'h0fce] = 8'hca;
s_mem_contents[14'h0fcf] = 8'he0;
s_mem_contents[14'h0fd0] = 8'hfa;
s_mem_contents[14'h0fd1] = 8'hb0;
s_mem_contents[14'h0fd2] = 8'hf6;
s_mem_contents[14'h0fd3] = 8'ha2;
s_mem_contents[14'h0fd4] = 8'h03;
s_mem_contents[14'h0fd5] = 8'ha0;
s_mem_contents[14'h0fd6] = 8'h00;
s_mem_contents[14'h0fd7] = 8'hb5;
s_mem_contents[14'h0fd8] = 8'h02;
s_mem_contents[14'h0fd9] = 8'hd5;
s_mem_contents[14'h0fda] = 8'h09;
s_mem_contents[14'h0fdb] = 8'hd0;
s_mem_contents[14'h0fdc] = 8'hfe;
s_mem_contents[14'h0fdd] = 8'h94;
s_mem_contents[14'h0fde] = 8'h02;
s_mem_contents[14'h0fdf] = 8'hbd;
s_mem_contents[14'h0fe0] = 8'h03;
s_mem_contents[14'h0fe1] = 8'h02;
s_mem_contents[14'h0fe2] = 8'hdd;
s_mem_contents[14'h0fe3] = 8'h17;
s_mem_contents[14'h0fe4] = 8'h02;
s_mem_contents[14'h0fe5] = 8'hd0;
s_mem_contents[14'h0fe6] = 8'hfe;
s_mem_contents[14'h0fe7] = 8'h8a;
s_mem_contents[14'h0fe8] = 8'h9d;
s_mem_contents[14'h0fe9] = 8'h03;
s_mem_contents[14'h0fea] = 8'h02;
s_mem_contents[14'h0feb] = 8'hca;
s_mem_contents[14'h0fec] = 8'h10;
s_mem_contents[14'h0fed] = 8'he9;
s_mem_contents[14'h0fee] = 8'had;
s_mem_contents[14'h0fef] = 8'h00;
s_mem_contents[14'h0ff0] = 8'h02;
s_mem_contents[14'h0ff1] = 8'hc9;
s_mem_contents[14'h0ff2] = 8'h12;
s_mem_contents[14'h0ff3] = 8'hd0;
s_mem_contents[14'h0ff4] = 8'hfe;
s_mem_contents[14'h0ff5] = 8'ha9;
s_mem_contents[14'h0ff6] = 8'h13;
s_mem_contents[14'h0ff7] = 8'h8d;
s_mem_contents[14'h0ff8] = 8'h00;
s_mem_contents[14'h0ff9] = 8'h02;
s_mem_contents[14'h0ffa] = 8'ha9;
s_mem_contents[14'h0ffb] = 8'h00;
s_mem_contents[14'h0ffc] = 8'h48;
s_mem_contents[14'h0ffd] = 8'h28;
s_mem_contents[14'h0ffe] = 8'ha6;
s_mem_contents[14'h0fff] = 8'h09;
s_mem_contents[14'h1000] = 8'h08;
s_mem_contents[14'h1001] = 8'h8a;
s_mem_contents[14'h1002] = 8'h49;
s_mem_contents[14'h1003] = 8'hc3;
s_mem_contents[14'h1004] = 8'haa;
s_mem_contents[14'h1005] = 8'h28;
s_mem_contents[14'h1006] = 8'h8e;
s_mem_contents[14'h1007] = 8'h03;
s_mem_contents[14'h1008] = 8'h02;
s_mem_contents[14'h1009] = 8'h08;
s_mem_contents[14'h100a] = 8'h49;
s_mem_contents[14'h100b] = 8'hc3;
s_mem_contents[14'h100c] = 8'haa;
s_mem_contents[14'h100d] = 8'he0;
s_mem_contents[14'h100e] = 8'hc3;
s_mem_contents[14'h100f] = 8'hd0;
s_mem_contents[14'h1010] = 8'hfe;
s_mem_contents[14'h1011] = 8'h68;
s_mem_contents[14'h1012] = 8'h49;
s_mem_contents[14'h1013] = 8'h30;
s_mem_contents[14'h1014] = 8'hcd;
s_mem_contents[14'h1015] = 8'h1c;
s_mem_contents[14'h1016] = 8'h02;
s_mem_contents[14'h1017] = 8'hd0;
s_mem_contents[14'h1018] = 8'hfe;
s_mem_contents[14'h1019] = 8'ha9;
s_mem_contents[14'h101a] = 8'h00;
s_mem_contents[14'h101b] = 8'h48;
s_mem_contents[14'h101c] = 8'h28;
s_mem_contents[14'h101d] = 8'ha6;
s_mem_contents[14'h101e] = 8'h0a;
s_mem_contents[14'h101f] = 8'h08;
s_mem_contents[14'h1020] = 8'h8a;
s_mem_contents[14'h1021] = 8'h49;
s_mem_contents[14'h1022] = 8'hc3;
s_mem_contents[14'h1023] = 8'haa;
s_mem_contents[14'h1024] = 8'h28;
s_mem_contents[14'h1025] = 8'h8e;
s_mem_contents[14'h1026] = 8'h04;
s_mem_contents[14'h1027] = 8'h02;
s_mem_contents[14'h1028] = 8'h08;
s_mem_contents[14'h1029] = 8'h49;
s_mem_contents[14'h102a] = 8'hc3;
s_mem_contents[14'h102b] = 8'haa;
s_mem_contents[14'h102c] = 8'he0;
s_mem_contents[14'h102d] = 8'h82;
s_mem_contents[14'h102e] = 8'hd0;
s_mem_contents[14'h102f] = 8'hfe;
s_mem_contents[14'h1030] = 8'h68;
s_mem_contents[14'h1031] = 8'h49;
s_mem_contents[14'h1032] = 8'h30;
s_mem_contents[14'h1033] = 8'hcd;
s_mem_contents[14'h1034] = 8'h1d;
s_mem_contents[14'h1035] = 8'h02;
s_mem_contents[14'h1036] = 8'hd0;
s_mem_contents[14'h1037] = 8'hfe;
s_mem_contents[14'h1038] = 8'ha9;
s_mem_contents[14'h1039] = 8'h00;
s_mem_contents[14'h103a] = 8'h48;
s_mem_contents[14'h103b] = 8'h28;
s_mem_contents[14'h103c] = 8'ha6;
s_mem_contents[14'h103d] = 8'h0b;
s_mem_contents[14'h103e] = 8'h08;
s_mem_contents[14'h103f] = 8'h8a;
s_mem_contents[14'h1040] = 8'h49;
s_mem_contents[14'h1041] = 8'hc3;
s_mem_contents[14'h1042] = 8'haa;
s_mem_contents[14'h1043] = 8'h28;
s_mem_contents[14'h1044] = 8'h8e;
s_mem_contents[14'h1045] = 8'h05;
s_mem_contents[14'h1046] = 8'h02;
s_mem_contents[14'h1047] = 8'h08;
s_mem_contents[14'h1048] = 8'h49;
s_mem_contents[14'h1049] = 8'hc3;
s_mem_contents[14'h104a] = 8'haa;
s_mem_contents[14'h104b] = 8'he0;
s_mem_contents[14'h104c] = 8'h41;
s_mem_contents[14'h104d] = 8'hd0;
s_mem_contents[14'h104e] = 8'hfe;
s_mem_contents[14'h104f] = 8'h68;
s_mem_contents[14'h1050] = 8'h49;
s_mem_contents[14'h1051] = 8'h30;
s_mem_contents[14'h1052] = 8'hcd;
s_mem_contents[14'h1053] = 8'h1e;
s_mem_contents[14'h1054] = 8'h02;
s_mem_contents[14'h1055] = 8'hd0;
s_mem_contents[14'h1056] = 8'hfe;
s_mem_contents[14'h1057] = 8'ha9;
s_mem_contents[14'h1058] = 8'h00;
s_mem_contents[14'h1059] = 8'h48;
s_mem_contents[14'h105a] = 8'h28;
s_mem_contents[14'h105b] = 8'ha6;
s_mem_contents[14'h105c] = 8'h0c;
s_mem_contents[14'h105d] = 8'h08;
s_mem_contents[14'h105e] = 8'h8a;
s_mem_contents[14'h105f] = 8'h49;
s_mem_contents[14'h1060] = 8'hc3;
s_mem_contents[14'h1061] = 8'haa;
s_mem_contents[14'h1062] = 8'h28;
s_mem_contents[14'h1063] = 8'h8e;
s_mem_contents[14'h1064] = 8'h06;
s_mem_contents[14'h1065] = 8'h02;
s_mem_contents[14'h1066] = 8'h08;
s_mem_contents[14'h1067] = 8'h49;
s_mem_contents[14'h1068] = 8'hc3;
s_mem_contents[14'h1069] = 8'haa;
s_mem_contents[14'h106a] = 8'he0;
s_mem_contents[14'h106b] = 8'h00;
s_mem_contents[14'h106c] = 8'hd0;
s_mem_contents[14'h106d] = 8'hfe;
s_mem_contents[14'h106e] = 8'h68;
s_mem_contents[14'h106f] = 8'h49;
s_mem_contents[14'h1070] = 8'h30;
s_mem_contents[14'h1071] = 8'hcd;
s_mem_contents[14'h1072] = 8'h1f;
s_mem_contents[14'h1073] = 8'h02;
s_mem_contents[14'h1074] = 8'hd0;
s_mem_contents[14'h1075] = 8'hfe;
s_mem_contents[14'h1076] = 8'ha9;
s_mem_contents[14'h1077] = 8'hff;
s_mem_contents[14'h1078] = 8'h48;
s_mem_contents[14'h1079] = 8'h28;
s_mem_contents[14'h107a] = 8'ha6;
s_mem_contents[14'h107b] = 8'h09;
s_mem_contents[14'h107c] = 8'h08;
s_mem_contents[14'h107d] = 8'h8a;
s_mem_contents[14'h107e] = 8'h49;
s_mem_contents[14'h107f] = 8'hc3;
s_mem_contents[14'h1080] = 8'haa;
s_mem_contents[14'h1081] = 8'h28;
s_mem_contents[14'h1082] = 8'h8e;
s_mem_contents[14'h1083] = 8'h03;
s_mem_contents[14'h1084] = 8'h02;
s_mem_contents[14'h1085] = 8'h08;
s_mem_contents[14'h1086] = 8'h49;
s_mem_contents[14'h1087] = 8'hc3;
s_mem_contents[14'h1088] = 8'haa;
s_mem_contents[14'h1089] = 8'he0;
s_mem_contents[14'h108a] = 8'hc3;
s_mem_contents[14'h108b] = 8'hd0;
s_mem_contents[14'h108c] = 8'hfe;
s_mem_contents[14'h108d] = 8'h68;
s_mem_contents[14'h108e] = 8'h49;
s_mem_contents[14'h108f] = 8'h7d;
s_mem_contents[14'h1090] = 8'hcd;
s_mem_contents[14'h1091] = 8'h1c;
s_mem_contents[14'h1092] = 8'h02;
s_mem_contents[14'h1093] = 8'hd0;
s_mem_contents[14'h1094] = 8'hfe;
s_mem_contents[14'h1095] = 8'ha9;
s_mem_contents[14'h1096] = 8'hff;
s_mem_contents[14'h1097] = 8'h48;
s_mem_contents[14'h1098] = 8'h28;
s_mem_contents[14'h1099] = 8'ha6;
s_mem_contents[14'h109a] = 8'h0a;
s_mem_contents[14'h109b] = 8'h08;
s_mem_contents[14'h109c] = 8'h8a;
s_mem_contents[14'h109d] = 8'h49;
s_mem_contents[14'h109e] = 8'hc3;
s_mem_contents[14'h109f] = 8'haa;
s_mem_contents[14'h10a0] = 8'h28;
s_mem_contents[14'h10a1] = 8'h8e;
s_mem_contents[14'h10a2] = 8'h04;
s_mem_contents[14'h10a3] = 8'h02;
s_mem_contents[14'h10a4] = 8'h08;
s_mem_contents[14'h10a5] = 8'h49;
s_mem_contents[14'h10a6] = 8'hc3;
s_mem_contents[14'h10a7] = 8'haa;
s_mem_contents[14'h10a8] = 8'he0;
s_mem_contents[14'h10a9] = 8'h82;
s_mem_contents[14'h10aa] = 8'hd0;
s_mem_contents[14'h10ab] = 8'hfe;
s_mem_contents[14'h10ac] = 8'h68;
s_mem_contents[14'h10ad] = 8'h49;
s_mem_contents[14'h10ae] = 8'h7d;
s_mem_contents[14'h10af] = 8'hcd;
s_mem_contents[14'h10b0] = 8'h1d;
s_mem_contents[14'h10b1] = 8'h02;
s_mem_contents[14'h10b2] = 8'hd0;
s_mem_contents[14'h10b3] = 8'hfe;
s_mem_contents[14'h10b4] = 8'ha9;
s_mem_contents[14'h10b5] = 8'hff;
s_mem_contents[14'h10b6] = 8'h48;
s_mem_contents[14'h10b7] = 8'h28;
s_mem_contents[14'h10b8] = 8'ha6;
s_mem_contents[14'h10b9] = 8'h0b;
s_mem_contents[14'h10ba] = 8'h08;
s_mem_contents[14'h10bb] = 8'h8a;
s_mem_contents[14'h10bc] = 8'h49;
s_mem_contents[14'h10bd] = 8'hc3;
s_mem_contents[14'h10be] = 8'haa;
s_mem_contents[14'h10bf] = 8'h28;
s_mem_contents[14'h10c0] = 8'h8e;
s_mem_contents[14'h10c1] = 8'h05;
s_mem_contents[14'h10c2] = 8'h02;
s_mem_contents[14'h10c3] = 8'h08;
s_mem_contents[14'h10c4] = 8'h49;
s_mem_contents[14'h10c5] = 8'hc3;
s_mem_contents[14'h10c6] = 8'haa;
s_mem_contents[14'h10c7] = 8'he0;
s_mem_contents[14'h10c8] = 8'h41;
s_mem_contents[14'h10c9] = 8'hd0;
s_mem_contents[14'h10ca] = 8'hfe;
s_mem_contents[14'h10cb] = 8'h68;
s_mem_contents[14'h10cc] = 8'h49;
s_mem_contents[14'h10cd] = 8'h7d;
s_mem_contents[14'h10ce] = 8'hcd;
s_mem_contents[14'h10cf] = 8'h1e;
s_mem_contents[14'h10d0] = 8'h02;
s_mem_contents[14'h10d1] = 8'hd0;
s_mem_contents[14'h10d2] = 8'hfe;
s_mem_contents[14'h10d3] = 8'ha9;
s_mem_contents[14'h10d4] = 8'hff;
s_mem_contents[14'h10d5] = 8'h48;
s_mem_contents[14'h10d6] = 8'h28;
s_mem_contents[14'h10d7] = 8'ha6;
s_mem_contents[14'h10d8] = 8'h0c;
s_mem_contents[14'h10d9] = 8'h08;
s_mem_contents[14'h10da] = 8'h8a;
s_mem_contents[14'h10db] = 8'h49;
s_mem_contents[14'h10dc] = 8'hc3;
s_mem_contents[14'h10dd] = 8'haa;
s_mem_contents[14'h10de] = 8'h28;
s_mem_contents[14'h10df] = 8'h8e;
s_mem_contents[14'h10e0] = 8'h06;
s_mem_contents[14'h10e1] = 8'h02;
s_mem_contents[14'h10e2] = 8'h08;
s_mem_contents[14'h10e3] = 8'h49;
s_mem_contents[14'h10e4] = 8'hc3;
s_mem_contents[14'h10e5] = 8'haa;
s_mem_contents[14'h10e6] = 8'he0;
s_mem_contents[14'h10e7] = 8'h00;
s_mem_contents[14'h10e8] = 8'hd0;
s_mem_contents[14'h10e9] = 8'hfe;
s_mem_contents[14'h10ea] = 8'h68;
s_mem_contents[14'h10eb] = 8'h49;
s_mem_contents[14'h10ec] = 8'h7d;
s_mem_contents[14'h10ed] = 8'hcd;
s_mem_contents[14'h10ee] = 8'h1f;
s_mem_contents[14'h10ef] = 8'h02;
s_mem_contents[14'h10f0] = 8'hd0;
s_mem_contents[14'h10f1] = 8'hfe;
s_mem_contents[14'h10f2] = 8'ha9;
s_mem_contents[14'h10f3] = 8'h00;
s_mem_contents[14'h10f4] = 8'h48;
s_mem_contents[14'h10f5] = 8'h28;
s_mem_contents[14'h10f6] = 8'hae;
s_mem_contents[14'h10f7] = 8'h17;
s_mem_contents[14'h10f8] = 8'h02;
s_mem_contents[14'h10f9] = 8'h08;
s_mem_contents[14'h10fa] = 8'h8a;
s_mem_contents[14'h10fb] = 8'h49;
s_mem_contents[14'h10fc] = 8'hc3;
s_mem_contents[14'h10fd] = 8'haa;
s_mem_contents[14'h10fe] = 8'h28;
s_mem_contents[14'h10ff] = 8'h86;
s_mem_contents[14'h1100] = 8'h02;
s_mem_contents[14'h1101] = 8'h08;
s_mem_contents[14'h1102] = 8'h49;
s_mem_contents[14'h1103] = 8'hc3;
s_mem_contents[14'h1104] = 8'hc5;
s_mem_contents[14'h1105] = 8'h09;
s_mem_contents[14'h1106] = 8'hd0;
s_mem_contents[14'h1107] = 8'hfe;
s_mem_contents[14'h1108] = 8'h68;
s_mem_contents[14'h1109] = 8'h49;
s_mem_contents[14'h110a] = 8'h30;
s_mem_contents[14'h110b] = 8'hcd;
s_mem_contents[14'h110c] = 8'h1c;
s_mem_contents[14'h110d] = 8'h02;
s_mem_contents[14'h110e] = 8'hd0;
s_mem_contents[14'h110f] = 8'hfe;
s_mem_contents[14'h1110] = 8'ha9;
s_mem_contents[14'h1111] = 8'h00;
s_mem_contents[14'h1112] = 8'h48;
s_mem_contents[14'h1113] = 8'h28;
s_mem_contents[14'h1114] = 8'hae;
s_mem_contents[14'h1115] = 8'h18;
s_mem_contents[14'h1116] = 8'h02;
s_mem_contents[14'h1117] = 8'h08;
s_mem_contents[14'h1118] = 8'h8a;
s_mem_contents[14'h1119] = 8'h49;
s_mem_contents[14'h111a] = 8'hc3;
s_mem_contents[14'h111b] = 8'haa;
s_mem_contents[14'h111c] = 8'h28;
s_mem_contents[14'h111d] = 8'h86;
s_mem_contents[14'h111e] = 8'h03;
s_mem_contents[14'h111f] = 8'h08;
s_mem_contents[14'h1120] = 8'h49;
s_mem_contents[14'h1121] = 8'hc3;
s_mem_contents[14'h1122] = 8'hc5;
s_mem_contents[14'h1123] = 8'h0a;
s_mem_contents[14'h1124] = 8'hd0;
s_mem_contents[14'h1125] = 8'hfe;
s_mem_contents[14'h1126] = 8'h68;
s_mem_contents[14'h1127] = 8'h49;
s_mem_contents[14'h1128] = 8'h30;
s_mem_contents[14'h1129] = 8'hcd;
s_mem_contents[14'h112a] = 8'h1d;
s_mem_contents[14'h112b] = 8'h02;
s_mem_contents[14'h112c] = 8'hd0;
s_mem_contents[14'h112d] = 8'hfe;
s_mem_contents[14'h112e] = 8'ha9;
s_mem_contents[14'h112f] = 8'h00;
s_mem_contents[14'h1130] = 8'h48;
s_mem_contents[14'h1131] = 8'h28;
s_mem_contents[14'h1132] = 8'hae;
s_mem_contents[14'h1133] = 8'h19;
s_mem_contents[14'h1134] = 8'h02;
s_mem_contents[14'h1135] = 8'h08;
s_mem_contents[14'h1136] = 8'h8a;
s_mem_contents[14'h1137] = 8'h49;
s_mem_contents[14'h1138] = 8'hc3;
s_mem_contents[14'h1139] = 8'haa;
s_mem_contents[14'h113a] = 8'h28;
s_mem_contents[14'h113b] = 8'h86;
s_mem_contents[14'h113c] = 8'h04;
s_mem_contents[14'h113d] = 8'h08;
s_mem_contents[14'h113e] = 8'h49;
s_mem_contents[14'h113f] = 8'hc3;
s_mem_contents[14'h1140] = 8'hc5;
s_mem_contents[14'h1141] = 8'h0b;
s_mem_contents[14'h1142] = 8'hd0;
s_mem_contents[14'h1143] = 8'hfe;
s_mem_contents[14'h1144] = 8'h68;
s_mem_contents[14'h1145] = 8'h49;
s_mem_contents[14'h1146] = 8'h30;
s_mem_contents[14'h1147] = 8'hcd;
s_mem_contents[14'h1148] = 8'h1e;
s_mem_contents[14'h1149] = 8'h02;
s_mem_contents[14'h114a] = 8'hd0;
s_mem_contents[14'h114b] = 8'hfe;
s_mem_contents[14'h114c] = 8'ha9;
s_mem_contents[14'h114d] = 8'h00;
s_mem_contents[14'h114e] = 8'h48;
s_mem_contents[14'h114f] = 8'h28;
s_mem_contents[14'h1150] = 8'hae;
s_mem_contents[14'h1151] = 8'h1a;
s_mem_contents[14'h1152] = 8'h02;
s_mem_contents[14'h1153] = 8'h08;
s_mem_contents[14'h1154] = 8'h8a;
s_mem_contents[14'h1155] = 8'h49;
s_mem_contents[14'h1156] = 8'hc3;
s_mem_contents[14'h1157] = 8'haa;
s_mem_contents[14'h1158] = 8'h28;
s_mem_contents[14'h1159] = 8'h86;
s_mem_contents[14'h115a] = 8'h05;
s_mem_contents[14'h115b] = 8'h08;
s_mem_contents[14'h115c] = 8'h49;
s_mem_contents[14'h115d] = 8'hc3;
s_mem_contents[14'h115e] = 8'hc5;
s_mem_contents[14'h115f] = 8'h0c;
s_mem_contents[14'h1160] = 8'hd0;
s_mem_contents[14'h1161] = 8'hfe;
s_mem_contents[14'h1162] = 8'h68;
s_mem_contents[14'h1163] = 8'h49;
s_mem_contents[14'h1164] = 8'h30;
s_mem_contents[14'h1165] = 8'hcd;
s_mem_contents[14'h1166] = 8'h1f;
s_mem_contents[14'h1167] = 8'h02;
s_mem_contents[14'h1168] = 8'hd0;
s_mem_contents[14'h1169] = 8'hfe;
s_mem_contents[14'h116a] = 8'ha9;
s_mem_contents[14'h116b] = 8'hff;
s_mem_contents[14'h116c] = 8'h48;
s_mem_contents[14'h116d] = 8'h28;
s_mem_contents[14'h116e] = 8'hae;
s_mem_contents[14'h116f] = 8'h17;
s_mem_contents[14'h1170] = 8'h02;
s_mem_contents[14'h1171] = 8'h08;
s_mem_contents[14'h1172] = 8'h8a;
s_mem_contents[14'h1173] = 8'h49;
s_mem_contents[14'h1174] = 8'hc3;
s_mem_contents[14'h1175] = 8'haa;
s_mem_contents[14'h1176] = 8'h28;
s_mem_contents[14'h1177] = 8'h86;
s_mem_contents[14'h1178] = 8'h02;
s_mem_contents[14'h1179] = 8'h08;
s_mem_contents[14'h117a] = 8'h49;
s_mem_contents[14'h117b] = 8'hc3;
s_mem_contents[14'h117c] = 8'haa;
s_mem_contents[14'h117d] = 8'he4;
s_mem_contents[14'h117e] = 8'h09;
s_mem_contents[14'h117f] = 8'hd0;
s_mem_contents[14'h1180] = 8'hfe;
s_mem_contents[14'h1181] = 8'h68;
s_mem_contents[14'h1182] = 8'h49;
s_mem_contents[14'h1183] = 8'h7d;
s_mem_contents[14'h1184] = 8'hcd;
s_mem_contents[14'h1185] = 8'h1c;
s_mem_contents[14'h1186] = 8'h02;
s_mem_contents[14'h1187] = 8'hd0;
s_mem_contents[14'h1188] = 8'hfe;
s_mem_contents[14'h1189] = 8'ha9;
s_mem_contents[14'h118a] = 8'hff;
s_mem_contents[14'h118b] = 8'h48;
s_mem_contents[14'h118c] = 8'h28;
s_mem_contents[14'h118d] = 8'hae;
s_mem_contents[14'h118e] = 8'h18;
s_mem_contents[14'h118f] = 8'h02;
s_mem_contents[14'h1190] = 8'h08;
s_mem_contents[14'h1191] = 8'h8a;
s_mem_contents[14'h1192] = 8'h49;
s_mem_contents[14'h1193] = 8'hc3;
s_mem_contents[14'h1194] = 8'haa;
s_mem_contents[14'h1195] = 8'h28;
s_mem_contents[14'h1196] = 8'h86;
s_mem_contents[14'h1197] = 8'h03;
s_mem_contents[14'h1198] = 8'h08;
s_mem_contents[14'h1199] = 8'h49;
s_mem_contents[14'h119a] = 8'hc3;
s_mem_contents[14'h119b] = 8'haa;
s_mem_contents[14'h119c] = 8'he4;
s_mem_contents[14'h119d] = 8'h0a;
s_mem_contents[14'h119e] = 8'hd0;
s_mem_contents[14'h119f] = 8'hfe;
s_mem_contents[14'h11a0] = 8'h68;
s_mem_contents[14'h11a1] = 8'h49;
s_mem_contents[14'h11a2] = 8'h7d;
s_mem_contents[14'h11a3] = 8'hcd;
s_mem_contents[14'h11a4] = 8'h1d;
s_mem_contents[14'h11a5] = 8'h02;
s_mem_contents[14'h11a6] = 8'hd0;
s_mem_contents[14'h11a7] = 8'hfe;
s_mem_contents[14'h11a8] = 8'ha9;
s_mem_contents[14'h11a9] = 8'hff;
s_mem_contents[14'h11aa] = 8'h48;
s_mem_contents[14'h11ab] = 8'h28;
s_mem_contents[14'h11ac] = 8'hae;
s_mem_contents[14'h11ad] = 8'h19;
s_mem_contents[14'h11ae] = 8'h02;
s_mem_contents[14'h11af] = 8'h08;
s_mem_contents[14'h11b0] = 8'h8a;
s_mem_contents[14'h11b1] = 8'h49;
s_mem_contents[14'h11b2] = 8'hc3;
s_mem_contents[14'h11b3] = 8'haa;
s_mem_contents[14'h11b4] = 8'h28;
s_mem_contents[14'h11b5] = 8'h86;
s_mem_contents[14'h11b6] = 8'h04;
s_mem_contents[14'h11b7] = 8'h08;
s_mem_contents[14'h11b8] = 8'h49;
s_mem_contents[14'h11b9] = 8'hc3;
s_mem_contents[14'h11ba] = 8'haa;
s_mem_contents[14'h11bb] = 8'he4;
s_mem_contents[14'h11bc] = 8'h0b;
s_mem_contents[14'h11bd] = 8'hd0;
s_mem_contents[14'h11be] = 8'hfe;
s_mem_contents[14'h11bf] = 8'h68;
s_mem_contents[14'h11c0] = 8'h49;
s_mem_contents[14'h11c1] = 8'h7d;
s_mem_contents[14'h11c2] = 8'hcd;
s_mem_contents[14'h11c3] = 8'h1e;
s_mem_contents[14'h11c4] = 8'h02;
s_mem_contents[14'h11c5] = 8'hd0;
s_mem_contents[14'h11c6] = 8'hfe;
s_mem_contents[14'h11c7] = 8'ha9;
s_mem_contents[14'h11c8] = 8'hff;
s_mem_contents[14'h11c9] = 8'h48;
s_mem_contents[14'h11ca] = 8'h28;
s_mem_contents[14'h11cb] = 8'hae;
s_mem_contents[14'h11cc] = 8'h1a;
s_mem_contents[14'h11cd] = 8'h02;
s_mem_contents[14'h11ce] = 8'h08;
s_mem_contents[14'h11cf] = 8'h8a;
s_mem_contents[14'h11d0] = 8'h49;
s_mem_contents[14'h11d1] = 8'hc3;
s_mem_contents[14'h11d2] = 8'haa;
s_mem_contents[14'h11d3] = 8'h28;
s_mem_contents[14'h11d4] = 8'h86;
s_mem_contents[14'h11d5] = 8'h05;
s_mem_contents[14'h11d6] = 8'h08;
s_mem_contents[14'h11d7] = 8'h49;
s_mem_contents[14'h11d8] = 8'hc3;
s_mem_contents[14'h11d9] = 8'haa;
s_mem_contents[14'h11da] = 8'he4;
s_mem_contents[14'h11db] = 8'h0c;
s_mem_contents[14'h11dc] = 8'hd0;
s_mem_contents[14'h11dd] = 8'hfe;
s_mem_contents[14'h11de] = 8'h68;
s_mem_contents[14'h11df] = 8'h49;
s_mem_contents[14'h11e0] = 8'h7d;
s_mem_contents[14'h11e1] = 8'hcd;
s_mem_contents[14'h11e2] = 8'h1f;
s_mem_contents[14'h11e3] = 8'h02;
s_mem_contents[14'h11e4] = 8'hd0;
s_mem_contents[14'h11e5] = 8'hfe;
s_mem_contents[14'h11e6] = 8'ha9;
s_mem_contents[14'h11e7] = 8'h00;
s_mem_contents[14'h11e8] = 8'h48;
s_mem_contents[14'h11e9] = 8'h28;
s_mem_contents[14'h11ea] = 8'ha2;
s_mem_contents[14'h11eb] = 8'hc3;
s_mem_contents[14'h11ec] = 8'h08;
s_mem_contents[14'h11ed] = 8'hec;
s_mem_contents[14'h11ee] = 8'h17;
s_mem_contents[14'h11ef] = 8'h02;
s_mem_contents[14'h11f0] = 8'hd0;
s_mem_contents[14'h11f1] = 8'hfe;
s_mem_contents[14'h11f2] = 8'h68;
s_mem_contents[14'h11f3] = 8'h49;
s_mem_contents[14'h11f4] = 8'h30;
s_mem_contents[14'h11f5] = 8'hcd;
s_mem_contents[14'h11f6] = 8'h1c;
s_mem_contents[14'h11f7] = 8'h02;
s_mem_contents[14'h11f8] = 8'hd0;
s_mem_contents[14'h11f9] = 8'hfe;
s_mem_contents[14'h11fa] = 8'ha9;
s_mem_contents[14'h11fb] = 8'h00;
s_mem_contents[14'h11fc] = 8'h48;
s_mem_contents[14'h11fd] = 8'h28;
s_mem_contents[14'h11fe] = 8'ha2;
s_mem_contents[14'h11ff] = 8'h82;
s_mem_contents[14'h1200] = 8'h08;
s_mem_contents[14'h1201] = 8'hec;
s_mem_contents[14'h1202] = 8'h18;
s_mem_contents[14'h1203] = 8'h02;
s_mem_contents[14'h1204] = 8'hd0;
s_mem_contents[14'h1205] = 8'hfe;
s_mem_contents[14'h1206] = 8'h68;
s_mem_contents[14'h1207] = 8'h49;
s_mem_contents[14'h1208] = 8'h30;
s_mem_contents[14'h1209] = 8'hcd;
s_mem_contents[14'h120a] = 8'h1d;
s_mem_contents[14'h120b] = 8'h02;
s_mem_contents[14'h120c] = 8'hd0;
s_mem_contents[14'h120d] = 8'hfe;
s_mem_contents[14'h120e] = 8'ha9;
s_mem_contents[14'h120f] = 8'h00;
s_mem_contents[14'h1210] = 8'h48;
s_mem_contents[14'h1211] = 8'h28;
s_mem_contents[14'h1212] = 8'ha2;
s_mem_contents[14'h1213] = 8'h41;
s_mem_contents[14'h1214] = 8'h08;
s_mem_contents[14'h1215] = 8'hec;
s_mem_contents[14'h1216] = 8'h19;
s_mem_contents[14'h1217] = 8'h02;
s_mem_contents[14'h1218] = 8'hd0;
s_mem_contents[14'h1219] = 8'hfe;
s_mem_contents[14'h121a] = 8'h68;
s_mem_contents[14'h121b] = 8'h49;
s_mem_contents[14'h121c] = 8'h30;
s_mem_contents[14'h121d] = 8'hcd;
s_mem_contents[14'h121e] = 8'h1e;
s_mem_contents[14'h121f] = 8'h02;
s_mem_contents[14'h1220] = 8'hd0;
s_mem_contents[14'h1221] = 8'hfe;
s_mem_contents[14'h1222] = 8'ha9;
s_mem_contents[14'h1223] = 8'h00;
s_mem_contents[14'h1224] = 8'h48;
s_mem_contents[14'h1225] = 8'h28;
s_mem_contents[14'h1226] = 8'ha2;
s_mem_contents[14'h1227] = 8'h00;
s_mem_contents[14'h1228] = 8'h08;
s_mem_contents[14'h1229] = 8'hec;
s_mem_contents[14'h122a] = 8'h1a;
s_mem_contents[14'h122b] = 8'h02;
s_mem_contents[14'h122c] = 8'hd0;
s_mem_contents[14'h122d] = 8'hfe;
s_mem_contents[14'h122e] = 8'h68;
s_mem_contents[14'h122f] = 8'h49;
s_mem_contents[14'h1230] = 8'h30;
s_mem_contents[14'h1231] = 8'hcd;
s_mem_contents[14'h1232] = 8'h1f;
s_mem_contents[14'h1233] = 8'h02;
s_mem_contents[14'h1234] = 8'hd0;
s_mem_contents[14'h1235] = 8'hfe;
s_mem_contents[14'h1236] = 8'ha9;
s_mem_contents[14'h1237] = 8'hff;
s_mem_contents[14'h1238] = 8'h48;
s_mem_contents[14'h1239] = 8'h28;
s_mem_contents[14'h123a] = 8'ha2;
s_mem_contents[14'h123b] = 8'hc3;
s_mem_contents[14'h123c] = 8'h08;
s_mem_contents[14'h123d] = 8'hec;
s_mem_contents[14'h123e] = 8'h17;
s_mem_contents[14'h123f] = 8'h02;
s_mem_contents[14'h1240] = 8'hd0;
s_mem_contents[14'h1241] = 8'hfe;
s_mem_contents[14'h1242] = 8'h68;
s_mem_contents[14'h1243] = 8'h49;
s_mem_contents[14'h1244] = 8'h7d;
s_mem_contents[14'h1245] = 8'hcd;
s_mem_contents[14'h1246] = 8'h1c;
s_mem_contents[14'h1247] = 8'h02;
s_mem_contents[14'h1248] = 8'hd0;
s_mem_contents[14'h1249] = 8'hfe;
s_mem_contents[14'h124a] = 8'ha9;
s_mem_contents[14'h124b] = 8'hff;
s_mem_contents[14'h124c] = 8'h48;
s_mem_contents[14'h124d] = 8'h28;
s_mem_contents[14'h124e] = 8'ha2;
s_mem_contents[14'h124f] = 8'h82;
s_mem_contents[14'h1250] = 8'h08;
s_mem_contents[14'h1251] = 8'hec;
s_mem_contents[14'h1252] = 8'h18;
s_mem_contents[14'h1253] = 8'h02;
s_mem_contents[14'h1254] = 8'hd0;
s_mem_contents[14'h1255] = 8'hfe;
s_mem_contents[14'h1256] = 8'h68;
s_mem_contents[14'h1257] = 8'h49;
s_mem_contents[14'h1258] = 8'h7d;
s_mem_contents[14'h1259] = 8'hcd;
s_mem_contents[14'h125a] = 8'h1d;
s_mem_contents[14'h125b] = 8'h02;
s_mem_contents[14'h125c] = 8'hd0;
s_mem_contents[14'h125d] = 8'hfe;
s_mem_contents[14'h125e] = 8'ha9;
s_mem_contents[14'h125f] = 8'hff;
s_mem_contents[14'h1260] = 8'h48;
s_mem_contents[14'h1261] = 8'h28;
s_mem_contents[14'h1262] = 8'ha2;
s_mem_contents[14'h1263] = 8'h41;
s_mem_contents[14'h1264] = 8'h08;
s_mem_contents[14'h1265] = 8'hec;
s_mem_contents[14'h1266] = 8'h19;
s_mem_contents[14'h1267] = 8'h02;
s_mem_contents[14'h1268] = 8'hd0;
s_mem_contents[14'h1269] = 8'hfe;
s_mem_contents[14'h126a] = 8'h68;
s_mem_contents[14'h126b] = 8'h49;
s_mem_contents[14'h126c] = 8'h7d;
s_mem_contents[14'h126d] = 8'hcd;
s_mem_contents[14'h126e] = 8'h1e;
s_mem_contents[14'h126f] = 8'h02;
s_mem_contents[14'h1270] = 8'hd0;
s_mem_contents[14'h1271] = 8'hfe;
s_mem_contents[14'h1272] = 8'ha9;
s_mem_contents[14'h1273] = 8'hff;
s_mem_contents[14'h1274] = 8'h48;
s_mem_contents[14'h1275] = 8'h28;
s_mem_contents[14'h1276] = 8'ha2;
s_mem_contents[14'h1277] = 8'h00;
s_mem_contents[14'h1278] = 8'h08;
s_mem_contents[14'h1279] = 8'hec;
s_mem_contents[14'h127a] = 8'h1a;
s_mem_contents[14'h127b] = 8'h02;
s_mem_contents[14'h127c] = 8'hd0;
s_mem_contents[14'h127d] = 8'hfe;
s_mem_contents[14'h127e] = 8'h68;
s_mem_contents[14'h127f] = 8'h49;
s_mem_contents[14'h1280] = 8'h7d;
s_mem_contents[14'h1281] = 8'hcd;
s_mem_contents[14'h1282] = 8'h1f;
s_mem_contents[14'h1283] = 8'h02;
s_mem_contents[14'h1284] = 8'hd0;
s_mem_contents[14'h1285] = 8'hfe;
s_mem_contents[14'h1286] = 8'ha2;
s_mem_contents[14'h1287] = 8'h00;
s_mem_contents[14'h1288] = 8'ha5;
s_mem_contents[14'h1289] = 8'h02;
s_mem_contents[14'h128a] = 8'h49;
s_mem_contents[14'h128b] = 8'hc3;
s_mem_contents[14'h128c] = 8'hc5;
s_mem_contents[14'h128d] = 8'h09;
s_mem_contents[14'h128e] = 8'hd0;
s_mem_contents[14'h128f] = 8'hfe;
s_mem_contents[14'h1290] = 8'h86;
s_mem_contents[14'h1291] = 8'h02;
s_mem_contents[14'h1292] = 8'had;
s_mem_contents[14'h1293] = 8'h03;
s_mem_contents[14'h1294] = 8'h02;
s_mem_contents[14'h1295] = 8'h49;
s_mem_contents[14'h1296] = 8'hc3;
s_mem_contents[14'h1297] = 8'hcd;
s_mem_contents[14'h1298] = 8'h17;
s_mem_contents[14'h1299] = 8'h02;
s_mem_contents[14'h129a] = 8'hd0;
s_mem_contents[14'h129b] = 8'hfe;
s_mem_contents[14'h129c] = 8'h8e;
s_mem_contents[14'h129d] = 8'h03;
s_mem_contents[14'h129e] = 8'h02;
s_mem_contents[14'h129f] = 8'ha5;
s_mem_contents[14'h12a0] = 8'h03;
s_mem_contents[14'h12a1] = 8'h49;
s_mem_contents[14'h12a2] = 8'hc3;
s_mem_contents[14'h12a3] = 8'hc5;
s_mem_contents[14'h12a4] = 8'h0a;
s_mem_contents[14'h12a5] = 8'hd0;
s_mem_contents[14'h12a6] = 8'hfe;
s_mem_contents[14'h12a7] = 8'h86;
s_mem_contents[14'h12a8] = 8'h03;
s_mem_contents[14'h12a9] = 8'had;
s_mem_contents[14'h12aa] = 8'h04;
s_mem_contents[14'h12ab] = 8'h02;
s_mem_contents[14'h12ac] = 8'h49;
s_mem_contents[14'h12ad] = 8'hc3;
s_mem_contents[14'h12ae] = 8'hcd;
s_mem_contents[14'h12af] = 8'h18;
s_mem_contents[14'h12b0] = 8'h02;
s_mem_contents[14'h12b1] = 8'hd0;
s_mem_contents[14'h12b2] = 8'hfe;
s_mem_contents[14'h12b3] = 8'h8e;
s_mem_contents[14'h12b4] = 8'h04;
s_mem_contents[14'h12b5] = 8'h02;
s_mem_contents[14'h12b6] = 8'ha5;
s_mem_contents[14'h12b7] = 8'h04;
s_mem_contents[14'h12b8] = 8'h49;
s_mem_contents[14'h12b9] = 8'hc3;
s_mem_contents[14'h12ba] = 8'hc5;
s_mem_contents[14'h12bb] = 8'h0b;
s_mem_contents[14'h12bc] = 8'hd0;
s_mem_contents[14'h12bd] = 8'hfe;
s_mem_contents[14'h12be] = 8'h86;
s_mem_contents[14'h12bf] = 8'h04;
s_mem_contents[14'h12c0] = 8'had;
s_mem_contents[14'h12c1] = 8'h05;
s_mem_contents[14'h12c2] = 8'h02;
s_mem_contents[14'h12c3] = 8'h49;
s_mem_contents[14'h12c4] = 8'hc3;
s_mem_contents[14'h12c5] = 8'hcd;
s_mem_contents[14'h12c6] = 8'h19;
s_mem_contents[14'h12c7] = 8'h02;
s_mem_contents[14'h12c8] = 8'hd0;
s_mem_contents[14'h12c9] = 8'hfe;
s_mem_contents[14'h12ca] = 8'h8e;
s_mem_contents[14'h12cb] = 8'h05;
s_mem_contents[14'h12cc] = 8'h02;
s_mem_contents[14'h12cd] = 8'ha5;
s_mem_contents[14'h12ce] = 8'h05;
s_mem_contents[14'h12cf] = 8'h49;
s_mem_contents[14'h12d0] = 8'hc3;
s_mem_contents[14'h12d1] = 8'hc5;
s_mem_contents[14'h12d2] = 8'h0c;
s_mem_contents[14'h12d3] = 8'hd0;
s_mem_contents[14'h12d4] = 8'hfe;
s_mem_contents[14'h12d5] = 8'h86;
s_mem_contents[14'h12d6] = 8'h05;
s_mem_contents[14'h12d7] = 8'had;
s_mem_contents[14'h12d8] = 8'h06;
s_mem_contents[14'h12d9] = 8'h02;
s_mem_contents[14'h12da] = 8'h49;
s_mem_contents[14'h12db] = 8'hc3;
s_mem_contents[14'h12dc] = 8'hcd;
s_mem_contents[14'h12dd] = 8'h1a;
s_mem_contents[14'h12de] = 8'h02;
s_mem_contents[14'h12df] = 8'hd0;
s_mem_contents[14'h12e0] = 8'hfe;
s_mem_contents[14'h12e1] = 8'h8e;
s_mem_contents[14'h12e2] = 8'h06;
s_mem_contents[14'h12e3] = 8'h02;
s_mem_contents[14'h12e4] = 8'had;
s_mem_contents[14'h12e5] = 8'h00;
s_mem_contents[14'h12e6] = 8'h02;
s_mem_contents[14'h12e7] = 8'hc9;
s_mem_contents[14'h12e8] = 8'h13;
s_mem_contents[14'h12e9] = 8'hd0;
s_mem_contents[14'h12ea] = 8'hfe;
s_mem_contents[14'h12eb] = 8'ha9;
s_mem_contents[14'h12ec] = 8'h14;
s_mem_contents[14'h12ed] = 8'h8d;
s_mem_contents[14'h12ee] = 8'h00;
s_mem_contents[14'h12ef] = 8'h02;
s_mem_contents[14'h12f0] = 8'ha9;
s_mem_contents[14'h12f1] = 8'h00;
s_mem_contents[14'h12f2] = 8'h48;
s_mem_contents[14'h12f3] = 8'h28;
s_mem_contents[14'h12f4] = 8'ha4;
s_mem_contents[14'h12f5] = 8'h09;
s_mem_contents[14'h12f6] = 8'h08;
s_mem_contents[14'h12f7] = 8'h98;
s_mem_contents[14'h12f8] = 8'h49;
s_mem_contents[14'h12f9] = 8'hc3;
s_mem_contents[14'h12fa] = 8'ha8;
s_mem_contents[14'h12fb] = 8'h28;
s_mem_contents[14'h12fc] = 8'h8c;
s_mem_contents[14'h12fd] = 8'h03;
s_mem_contents[14'h12fe] = 8'h02;
s_mem_contents[14'h12ff] = 8'h08;
s_mem_contents[14'h1300] = 8'h49;
s_mem_contents[14'h1301] = 8'hc3;
s_mem_contents[14'h1302] = 8'ha8;
s_mem_contents[14'h1303] = 8'hc0;
s_mem_contents[14'h1304] = 8'hc3;
s_mem_contents[14'h1305] = 8'hd0;
s_mem_contents[14'h1306] = 8'hfe;
s_mem_contents[14'h1307] = 8'h68;
s_mem_contents[14'h1308] = 8'h49;
s_mem_contents[14'h1309] = 8'h30;
s_mem_contents[14'h130a] = 8'hcd;
s_mem_contents[14'h130b] = 8'h1c;
s_mem_contents[14'h130c] = 8'h02;
s_mem_contents[14'h130d] = 8'hd0;
s_mem_contents[14'h130e] = 8'hfe;
s_mem_contents[14'h130f] = 8'ha9;
s_mem_contents[14'h1310] = 8'h00;
s_mem_contents[14'h1311] = 8'h48;
s_mem_contents[14'h1312] = 8'h28;
s_mem_contents[14'h1313] = 8'ha4;
s_mem_contents[14'h1314] = 8'h0a;
s_mem_contents[14'h1315] = 8'h08;
s_mem_contents[14'h1316] = 8'h98;
s_mem_contents[14'h1317] = 8'h49;
s_mem_contents[14'h1318] = 8'hc3;
s_mem_contents[14'h1319] = 8'ha8;
s_mem_contents[14'h131a] = 8'h28;
s_mem_contents[14'h131b] = 8'h8c;
s_mem_contents[14'h131c] = 8'h04;
s_mem_contents[14'h131d] = 8'h02;
s_mem_contents[14'h131e] = 8'h08;
s_mem_contents[14'h131f] = 8'h49;
s_mem_contents[14'h1320] = 8'hc3;
s_mem_contents[14'h1321] = 8'ha8;
s_mem_contents[14'h1322] = 8'hc0;
s_mem_contents[14'h1323] = 8'h82;
s_mem_contents[14'h1324] = 8'hd0;
s_mem_contents[14'h1325] = 8'hfe;
s_mem_contents[14'h1326] = 8'h68;
s_mem_contents[14'h1327] = 8'h49;
s_mem_contents[14'h1328] = 8'h30;
s_mem_contents[14'h1329] = 8'hcd;
s_mem_contents[14'h132a] = 8'h1d;
s_mem_contents[14'h132b] = 8'h02;
s_mem_contents[14'h132c] = 8'hd0;
s_mem_contents[14'h132d] = 8'hfe;
s_mem_contents[14'h132e] = 8'ha9;
s_mem_contents[14'h132f] = 8'h00;
s_mem_contents[14'h1330] = 8'h48;
s_mem_contents[14'h1331] = 8'h28;
s_mem_contents[14'h1332] = 8'ha4;
s_mem_contents[14'h1333] = 8'h0b;
s_mem_contents[14'h1334] = 8'h08;
s_mem_contents[14'h1335] = 8'h98;
s_mem_contents[14'h1336] = 8'h49;
s_mem_contents[14'h1337] = 8'hc3;
s_mem_contents[14'h1338] = 8'ha8;
s_mem_contents[14'h1339] = 8'h28;
s_mem_contents[14'h133a] = 8'h8c;
s_mem_contents[14'h133b] = 8'h05;
s_mem_contents[14'h133c] = 8'h02;
s_mem_contents[14'h133d] = 8'h08;
s_mem_contents[14'h133e] = 8'h49;
s_mem_contents[14'h133f] = 8'hc3;
s_mem_contents[14'h1340] = 8'ha8;
s_mem_contents[14'h1341] = 8'hc0;
s_mem_contents[14'h1342] = 8'h41;
s_mem_contents[14'h1343] = 8'hd0;
s_mem_contents[14'h1344] = 8'hfe;
s_mem_contents[14'h1345] = 8'h68;
s_mem_contents[14'h1346] = 8'h49;
s_mem_contents[14'h1347] = 8'h30;
s_mem_contents[14'h1348] = 8'hcd;
s_mem_contents[14'h1349] = 8'h1e;
s_mem_contents[14'h134a] = 8'h02;
s_mem_contents[14'h134b] = 8'hd0;
s_mem_contents[14'h134c] = 8'hfe;
s_mem_contents[14'h134d] = 8'ha9;
s_mem_contents[14'h134e] = 8'h00;
s_mem_contents[14'h134f] = 8'h48;
s_mem_contents[14'h1350] = 8'h28;
s_mem_contents[14'h1351] = 8'ha4;
s_mem_contents[14'h1352] = 8'h0c;
s_mem_contents[14'h1353] = 8'h08;
s_mem_contents[14'h1354] = 8'h98;
s_mem_contents[14'h1355] = 8'h49;
s_mem_contents[14'h1356] = 8'hc3;
s_mem_contents[14'h1357] = 8'ha8;
s_mem_contents[14'h1358] = 8'h28;
s_mem_contents[14'h1359] = 8'h8c;
s_mem_contents[14'h135a] = 8'h06;
s_mem_contents[14'h135b] = 8'h02;
s_mem_contents[14'h135c] = 8'h08;
s_mem_contents[14'h135d] = 8'h49;
s_mem_contents[14'h135e] = 8'hc3;
s_mem_contents[14'h135f] = 8'ha8;
s_mem_contents[14'h1360] = 8'hc0;
s_mem_contents[14'h1361] = 8'h00;
s_mem_contents[14'h1362] = 8'hd0;
s_mem_contents[14'h1363] = 8'hfe;
s_mem_contents[14'h1364] = 8'h68;
s_mem_contents[14'h1365] = 8'h49;
s_mem_contents[14'h1366] = 8'h30;
s_mem_contents[14'h1367] = 8'hcd;
s_mem_contents[14'h1368] = 8'h1f;
s_mem_contents[14'h1369] = 8'h02;
s_mem_contents[14'h136a] = 8'hd0;
s_mem_contents[14'h136b] = 8'hfe;
s_mem_contents[14'h136c] = 8'ha9;
s_mem_contents[14'h136d] = 8'hff;
s_mem_contents[14'h136e] = 8'h48;
s_mem_contents[14'h136f] = 8'h28;
s_mem_contents[14'h1370] = 8'ha4;
s_mem_contents[14'h1371] = 8'h09;
s_mem_contents[14'h1372] = 8'h08;
s_mem_contents[14'h1373] = 8'h98;
s_mem_contents[14'h1374] = 8'h49;
s_mem_contents[14'h1375] = 8'hc3;
s_mem_contents[14'h1376] = 8'ha8;
s_mem_contents[14'h1377] = 8'h28;
s_mem_contents[14'h1378] = 8'h8c;
s_mem_contents[14'h1379] = 8'h03;
s_mem_contents[14'h137a] = 8'h02;
s_mem_contents[14'h137b] = 8'h08;
s_mem_contents[14'h137c] = 8'h49;
s_mem_contents[14'h137d] = 8'hc3;
s_mem_contents[14'h137e] = 8'ha8;
s_mem_contents[14'h137f] = 8'hc0;
s_mem_contents[14'h1380] = 8'hc3;
s_mem_contents[14'h1381] = 8'hd0;
s_mem_contents[14'h1382] = 8'hfe;
s_mem_contents[14'h1383] = 8'h68;
s_mem_contents[14'h1384] = 8'h49;
s_mem_contents[14'h1385] = 8'h7d;
s_mem_contents[14'h1386] = 8'hcd;
s_mem_contents[14'h1387] = 8'h1c;
s_mem_contents[14'h1388] = 8'h02;
s_mem_contents[14'h1389] = 8'hd0;
s_mem_contents[14'h138a] = 8'hfe;
s_mem_contents[14'h138b] = 8'ha9;
s_mem_contents[14'h138c] = 8'hff;
s_mem_contents[14'h138d] = 8'h48;
s_mem_contents[14'h138e] = 8'h28;
s_mem_contents[14'h138f] = 8'ha4;
s_mem_contents[14'h1390] = 8'h0a;
s_mem_contents[14'h1391] = 8'h08;
s_mem_contents[14'h1392] = 8'h98;
s_mem_contents[14'h1393] = 8'h49;
s_mem_contents[14'h1394] = 8'hc3;
s_mem_contents[14'h1395] = 8'ha8;
s_mem_contents[14'h1396] = 8'h28;
s_mem_contents[14'h1397] = 8'h8c;
s_mem_contents[14'h1398] = 8'h04;
s_mem_contents[14'h1399] = 8'h02;
s_mem_contents[14'h139a] = 8'h08;
s_mem_contents[14'h139b] = 8'h49;
s_mem_contents[14'h139c] = 8'hc3;
s_mem_contents[14'h139d] = 8'ha8;
s_mem_contents[14'h139e] = 8'hc0;
s_mem_contents[14'h139f] = 8'h82;
s_mem_contents[14'h13a0] = 8'hd0;
s_mem_contents[14'h13a1] = 8'hfe;
s_mem_contents[14'h13a2] = 8'h68;
s_mem_contents[14'h13a3] = 8'h49;
s_mem_contents[14'h13a4] = 8'h7d;
s_mem_contents[14'h13a5] = 8'hcd;
s_mem_contents[14'h13a6] = 8'h1d;
s_mem_contents[14'h13a7] = 8'h02;
s_mem_contents[14'h13a8] = 8'hd0;
s_mem_contents[14'h13a9] = 8'hfe;
s_mem_contents[14'h13aa] = 8'ha9;
s_mem_contents[14'h13ab] = 8'hff;
s_mem_contents[14'h13ac] = 8'h48;
s_mem_contents[14'h13ad] = 8'h28;
s_mem_contents[14'h13ae] = 8'ha4;
s_mem_contents[14'h13af] = 8'h0b;
s_mem_contents[14'h13b0] = 8'h08;
s_mem_contents[14'h13b1] = 8'h98;
s_mem_contents[14'h13b2] = 8'h49;
s_mem_contents[14'h13b3] = 8'hc3;
s_mem_contents[14'h13b4] = 8'ha8;
s_mem_contents[14'h13b5] = 8'h28;
s_mem_contents[14'h13b6] = 8'h8c;
s_mem_contents[14'h13b7] = 8'h05;
s_mem_contents[14'h13b8] = 8'h02;
s_mem_contents[14'h13b9] = 8'h08;
s_mem_contents[14'h13ba] = 8'h49;
s_mem_contents[14'h13bb] = 8'hc3;
s_mem_contents[14'h13bc] = 8'ha8;
s_mem_contents[14'h13bd] = 8'hc0;
s_mem_contents[14'h13be] = 8'h41;
s_mem_contents[14'h13bf] = 8'hd0;
s_mem_contents[14'h13c0] = 8'hfe;
s_mem_contents[14'h13c1] = 8'h68;
s_mem_contents[14'h13c2] = 8'h49;
s_mem_contents[14'h13c3] = 8'h7d;
s_mem_contents[14'h13c4] = 8'hcd;
s_mem_contents[14'h13c5] = 8'h1e;
s_mem_contents[14'h13c6] = 8'h02;
s_mem_contents[14'h13c7] = 8'hd0;
s_mem_contents[14'h13c8] = 8'hfe;
s_mem_contents[14'h13c9] = 8'ha9;
s_mem_contents[14'h13ca] = 8'hff;
s_mem_contents[14'h13cb] = 8'h48;
s_mem_contents[14'h13cc] = 8'h28;
s_mem_contents[14'h13cd] = 8'ha4;
s_mem_contents[14'h13ce] = 8'h0c;
s_mem_contents[14'h13cf] = 8'h08;
s_mem_contents[14'h13d0] = 8'h98;
s_mem_contents[14'h13d1] = 8'h49;
s_mem_contents[14'h13d2] = 8'hc3;
s_mem_contents[14'h13d3] = 8'ha8;
s_mem_contents[14'h13d4] = 8'h28;
s_mem_contents[14'h13d5] = 8'h8c;
s_mem_contents[14'h13d6] = 8'h06;
s_mem_contents[14'h13d7] = 8'h02;
s_mem_contents[14'h13d8] = 8'h08;
s_mem_contents[14'h13d9] = 8'h49;
s_mem_contents[14'h13da] = 8'hc3;
s_mem_contents[14'h13db] = 8'ha8;
s_mem_contents[14'h13dc] = 8'hc0;
s_mem_contents[14'h13dd] = 8'h00;
s_mem_contents[14'h13de] = 8'hd0;
s_mem_contents[14'h13df] = 8'hfe;
s_mem_contents[14'h13e0] = 8'h68;
s_mem_contents[14'h13e1] = 8'h49;
s_mem_contents[14'h13e2] = 8'h7d;
s_mem_contents[14'h13e3] = 8'hcd;
s_mem_contents[14'h13e4] = 8'h1f;
s_mem_contents[14'h13e5] = 8'h02;
s_mem_contents[14'h13e6] = 8'hd0;
s_mem_contents[14'h13e7] = 8'hfe;
s_mem_contents[14'h13e8] = 8'ha9;
s_mem_contents[14'h13e9] = 8'h00;
s_mem_contents[14'h13ea] = 8'h48;
s_mem_contents[14'h13eb] = 8'h28;
s_mem_contents[14'h13ec] = 8'hac;
s_mem_contents[14'h13ed] = 8'h17;
s_mem_contents[14'h13ee] = 8'h02;
s_mem_contents[14'h13ef] = 8'h08;
s_mem_contents[14'h13f0] = 8'h98;
s_mem_contents[14'h13f1] = 8'h49;
s_mem_contents[14'h13f2] = 8'hc3;
s_mem_contents[14'h13f3] = 8'ha8;
s_mem_contents[14'h13f4] = 8'h28;
s_mem_contents[14'h13f5] = 8'h84;
s_mem_contents[14'h13f6] = 8'h02;
s_mem_contents[14'h13f7] = 8'h08;
s_mem_contents[14'h13f8] = 8'h49;
s_mem_contents[14'h13f9] = 8'hc3;
s_mem_contents[14'h13fa] = 8'ha8;
s_mem_contents[14'h13fb] = 8'hc4;
s_mem_contents[14'h13fc] = 8'h09;
s_mem_contents[14'h13fd] = 8'hd0;
s_mem_contents[14'h13fe] = 8'hfe;
s_mem_contents[14'h13ff] = 8'h68;
s_mem_contents[14'h1400] = 8'h49;
s_mem_contents[14'h1401] = 8'h30;
s_mem_contents[14'h1402] = 8'hcd;
s_mem_contents[14'h1403] = 8'h1c;
s_mem_contents[14'h1404] = 8'h02;
s_mem_contents[14'h1405] = 8'hd0;
s_mem_contents[14'h1406] = 8'hfe;
s_mem_contents[14'h1407] = 8'ha9;
s_mem_contents[14'h1408] = 8'h00;
s_mem_contents[14'h1409] = 8'h48;
s_mem_contents[14'h140a] = 8'h28;
s_mem_contents[14'h140b] = 8'hac;
s_mem_contents[14'h140c] = 8'h18;
s_mem_contents[14'h140d] = 8'h02;
s_mem_contents[14'h140e] = 8'h08;
s_mem_contents[14'h140f] = 8'h98;
s_mem_contents[14'h1410] = 8'h49;
s_mem_contents[14'h1411] = 8'hc3;
s_mem_contents[14'h1412] = 8'ha8;
s_mem_contents[14'h1413] = 8'h28;
s_mem_contents[14'h1414] = 8'h84;
s_mem_contents[14'h1415] = 8'h03;
s_mem_contents[14'h1416] = 8'h08;
s_mem_contents[14'h1417] = 8'h49;
s_mem_contents[14'h1418] = 8'hc3;
s_mem_contents[14'h1419] = 8'ha8;
s_mem_contents[14'h141a] = 8'hc4;
s_mem_contents[14'h141b] = 8'h0a;
s_mem_contents[14'h141c] = 8'hd0;
s_mem_contents[14'h141d] = 8'hfe;
s_mem_contents[14'h141e] = 8'h68;
s_mem_contents[14'h141f] = 8'h49;
s_mem_contents[14'h1420] = 8'h30;
s_mem_contents[14'h1421] = 8'hcd;
s_mem_contents[14'h1422] = 8'h1d;
s_mem_contents[14'h1423] = 8'h02;
s_mem_contents[14'h1424] = 8'hd0;
s_mem_contents[14'h1425] = 8'hfe;
s_mem_contents[14'h1426] = 8'ha9;
s_mem_contents[14'h1427] = 8'h00;
s_mem_contents[14'h1428] = 8'h48;
s_mem_contents[14'h1429] = 8'h28;
s_mem_contents[14'h142a] = 8'hac;
s_mem_contents[14'h142b] = 8'h19;
s_mem_contents[14'h142c] = 8'h02;
s_mem_contents[14'h142d] = 8'h08;
s_mem_contents[14'h142e] = 8'h98;
s_mem_contents[14'h142f] = 8'h49;
s_mem_contents[14'h1430] = 8'hc3;
s_mem_contents[14'h1431] = 8'ha8;
s_mem_contents[14'h1432] = 8'h28;
s_mem_contents[14'h1433] = 8'h84;
s_mem_contents[14'h1434] = 8'h04;
s_mem_contents[14'h1435] = 8'h08;
s_mem_contents[14'h1436] = 8'h49;
s_mem_contents[14'h1437] = 8'hc3;
s_mem_contents[14'h1438] = 8'ha8;
s_mem_contents[14'h1439] = 8'hc4;
s_mem_contents[14'h143a] = 8'h0b;
s_mem_contents[14'h143b] = 8'hd0;
s_mem_contents[14'h143c] = 8'hfe;
s_mem_contents[14'h143d] = 8'h68;
s_mem_contents[14'h143e] = 8'h49;
s_mem_contents[14'h143f] = 8'h30;
s_mem_contents[14'h1440] = 8'hcd;
s_mem_contents[14'h1441] = 8'h1e;
s_mem_contents[14'h1442] = 8'h02;
s_mem_contents[14'h1443] = 8'hd0;
s_mem_contents[14'h1444] = 8'hfe;
s_mem_contents[14'h1445] = 8'ha9;
s_mem_contents[14'h1446] = 8'h00;
s_mem_contents[14'h1447] = 8'h48;
s_mem_contents[14'h1448] = 8'h28;
s_mem_contents[14'h1449] = 8'hac;
s_mem_contents[14'h144a] = 8'h1a;
s_mem_contents[14'h144b] = 8'h02;
s_mem_contents[14'h144c] = 8'h08;
s_mem_contents[14'h144d] = 8'h98;
s_mem_contents[14'h144e] = 8'h49;
s_mem_contents[14'h144f] = 8'hc3;
s_mem_contents[14'h1450] = 8'ha8;
s_mem_contents[14'h1451] = 8'h28;
s_mem_contents[14'h1452] = 8'h84;
s_mem_contents[14'h1453] = 8'h05;
s_mem_contents[14'h1454] = 8'h08;
s_mem_contents[14'h1455] = 8'h49;
s_mem_contents[14'h1456] = 8'hc3;
s_mem_contents[14'h1457] = 8'ha8;
s_mem_contents[14'h1458] = 8'hc4;
s_mem_contents[14'h1459] = 8'h0c;
s_mem_contents[14'h145a] = 8'hd0;
s_mem_contents[14'h145b] = 8'hfe;
s_mem_contents[14'h145c] = 8'h68;
s_mem_contents[14'h145d] = 8'h49;
s_mem_contents[14'h145e] = 8'h30;
s_mem_contents[14'h145f] = 8'hcd;
s_mem_contents[14'h1460] = 8'h1f;
s_mem_contents[14'h1461] = 8'h02;
s_mem_contents[14'h1462] = 8'hd0;
s_mem_contents[14'h1463] = 8'hfe;
s_mem_contents[14'h1464] = 8'ha9;
s_mem_contents[14'h1465] = 8'hff;
s_mem_contents[14'h1466] = 8'h48;
s_mem_contents[14'h1467] = 8'h28;
s_mem_contents[14'h1468] = 8'hac;
s_mem_contents[14'h1469] = 8'h17;
s_mem_contents[14'h146a] = 8'h02;
s_mem_contents[14'h146b] = 8'h08;
s_mem_contents[14'h146c] = 8'h98;
s_mem_contents[14'h146d] = 8'h49;
s_mem_contents[14'h146e] = 8'hc3;
s_mem_contents[14'h146f] = 8'ha8;
s_mem_contents[14'h1470] = 8'h28;
s_mem_contents[14'h1471] = 8'h84;
s_mem_contents[14'h1472] = 8'h02;
s_mem_contents[14'h1473] = 8'h08;
s_mem_contents[14'h1474] = 8'h49;
s_mem_contents[14'h1475] = 8'hc3;
s_mem_contents[14'h1476] = 8'ha8;
s_mem_contents[14'h1477] = 8'hc5;
s_mem_contents[14'h1478] = 8'h09;
s_mem_contents[14'h1479] = 8'hd0;
s_mem_contents[14'h147a] = 8'hfe;
s_mem_contents[14'h147b] = 8'h68;
s_mem_contents[14'h147c] = 8'h49;
s_mem_contents[14'h147d] = 8'h7d;
s_mem_contents[14'h147e] = 8'hcd;
s_mem_contents[14'h147f] = 8'h1c;
s_mem_contents[14'h1480] = 8'h02;
s_mem_contents[14'h1481] = 8'hd0;
s_mem_contents[14'h1482] = 8'hfe;
s_mem_contents[14'h1483] = 8'ha9;
s_mem_contents[14'h1484] = 8'hff;
s_mem_contents[14'h1485] = 8'h48;
s_mem_contents[14'h1486] = 8'h28;
s_mem_contents[14'h1487] = 8'hac;
s_mem_contents[14'h1488] = 8'h18;
s_mem_contents[14'h1489] = 8'h02;
s_mem_contents[14'h148a] = 8'h08;
s_mem_contents[14'h148b] = 8'h98;
s_mem_contents[14'h148c] = 8'h49;
s_mem_contents[14'h148d] = 8'hc3;
s_mem_contents[14'h148e] = 8'ha8;
s_mem_contents[14'h148f] = 8'h28;
s_mem_contents[14'h1490] = 8'h84;
s_mem_contents[14'h1491] = 8'h03;
s_mem_contents[14'h1492] = 8'h08;
s_mem_contents[14'h1493] = 8'h49;
s_mem_contents[14'h1494] = 8'hc3;
s_mem_contents[14'h1495] = 8'ha8;
s_mem_contents[14'h1496] = 8'hc5;
s_mem_contents[14'h1497] = 8'h0a;
s_mem_contents[14'h1498] = 8'hd0;
s_mem_contents[14'h1499] = 8'hfe;
s_mem_contents[14'h149a] = 8'h68;
s_mem_contents[14'h149b] = 8'h49;
s_mem_contents[14'h149c] = 8'h7d;
s_mem_contents[14'h149d] = 8'hcd;
s_mem_contents[14'h149e] = 8'h1d;
s_mem_contents[14'h149f] = 8'h02;
s_mem_contents[14'h14a0] = 8'hd0;
s_mem_contents[14'h14a1] = 8'hfe;
s_mem_contents[14'h14a2] = 8'ha9;
s_mem_contents[14'h14a3] = 8'hff;
s_mem_contents[14'h14a4] = 8'h48;
s_mem_contents[14'h14a5] = 8'h28;
s_mem_contents[14'h14a6] = 8'hac;
s_mem_contents[14'h14a7] = 8'h19;
s_mem_contents[14'h14a8] = 8'h02;
s_mem_contents[14'h14a9] = 8'h08;
s_mem_contents[14'h14aa] = 8'h98;
s_mem_contents[14'h14ab] = 8'h49;
s_mem_contents[14'h14ac] = 8'hc3;
s_mem_contents[14'h14ad] = 8'ha8;
s_mem_contents[14'h14ae] = 8'h28;
s_mem_contents[14'h14af] = 8'h84;
s_mem_contents[14'h14b0] = 8'h04;
s_mem_contents[14'h14b1] = 8'h08;
s_mem_contents[14'h14b2] = 8'h49;
s_mem_contents[14'h14b3] = 8'hc3;
s_mem_contents[14'h14b4] = 8'ha8;
s_mem_contents[14'h14b5] = 8'hc5;
s_mem_contents[14'h14b6] = 8'h0b;
s_mem_contents[14'h14b7] = 8'hd0;
s_mem_contents[14'h14b8] = 8'hfe;
s_mem_contents[14'h14b9] = 8'h68;
s_mem_contents[14'h14ba] = 8'h49;
s_mem_contents[14'h14bb] = 8'h7d;
s_mem_contents[14'h14bc] = 8'hcd;
s_mem_contents[14'h14bd] = 8'h1e;
s_mem_contents[14'h14be] = 8'h02;
s_mem_contents[14'h14bf] = 8'hd0;
s_mem_contents[14'h14c0] = 8'hfe;
s_mem_contents[14'h14c1] = 8'ha9;
s_mem_contents[14'h14c2] = 8'hff;
s_mem_contents[14'h14c3] = 8'h48;
s_mem_contents[14'h14c4] = 8'h28;
s_mem_contents[14'h14c5] = 8'hac;
s_mem_contents[14'h14c6] = 8'h1a;
s_mem_contents[14'h14c7] = 8'h02;
s_mem_contents[14'h14c8] = 8'h08;
s_mem_contents[14'h14c9] = 8'h98;
s_mem_contents[14'h14ca] = 8'h49;
s_mem_contents[14'h14cb] = 8'hc3;
s_mem_contents[14'h14cc] = 8'ha8;
s_mem_contents[14'h14cd] = 8'h28;
s_mem_contents[14'h14ce] = 8'h84;
s_mem_contents[14'h14cf] = 8'h05;
s_mem_contents[14'h14d0] = 8'h08;
s_mem_contents[14'h14d1] = 8'h49;
s_mem_contents[14'h14d2] = 8'hc3;
s_mem_contents[14'h14d3] = 8'ha8;
s_mem_contents[14'h14d4] = 8'hc5;
s_mem_contents[14'h14d5] = 8'h0c;
s_mem_contents[14'h14d6] = 8'hd0;
s_mem_contents[14'h14d7] = 8'hfe;
s_mem_contents[14'h14d8] = 8'h68;
s_mem_contents[14'h14d9] = 8'h49;
s_mem_contents[14'h14da] = 8'h7d;
s_mem_contents[14'h14db] = 8'hcd;
s_mem_contents[14'h14dc] = 8'h1f;
s_mem_contents[14'h14dd] = 8'h02;
s_mem_contents[14'h14de] = 8'hd0;
s_mem_contents[14'h14df] = 8'hfe;
s_mem_contents[14'h14e0] = 8'ha9;
s_mem_contents[14'h14e1] = 8'h00;
s_mem_contents[14'h14e2] = 8'h48;
s_mem_contents[14'h14e3] = 8'h28;
s_mem_contents[14'h14e4] = 8'ha0;
s_mem_contents[14'h14e5] = 8'hc3;
s_mem_contents[14'h14e6] = 8'h08;
s_mem_contents[14'h14e7] = 8'hcc;
s_mem_contents[14'h14e8] = 8'h17;
s_mem_contents[14'h14e9] = 8'h02;
s_mem_contents[14'h14ea] = 8'hd0;
s_mem_contents[14'h14eb] = 8'hfe;
s_mem_contents[14'h14ec] = 8'h68;
s_mem_contents[14'h14ed] = 8'h49;
s_mem_contents[14'h14ee] = 8'h30;
s_mem_contents[14'h14ef] = 8'hcd;
s_mem_contents[14'h14f0] = 8'h1c;
s_mem_contents[14'h14f1] = 8'h02;
s_mem_contents[14'h14f2] = 8'hd0;
s_mem_contents[14'h14f3] = 8'hfe;
s_mem_contents[14'h14f4] = 8'ha9;
s_mem_contents[14'h14f5] = 8'h00;
s_mem_contents[14'h14f6] = 8'h48;
s_mem_contents[14'h14f7] = 8'h28;
s_mem_contents[14'h14f8] = 8'ha0;
s_mem_contents[14'h14f9] = 8'h82;
s_mem_contents[14'h14fa] = 8'h08;
s_mem_contents[14'h14fb] = 8'hcc;
s_mem_contents[14'h14fc] = 8'h18;
s_mem_contents[14'h14fd] = 8'h02;
s_mem_contents[14'h14fe] = 8'hd0;
s_mem_contents[14'h14ff] = 8'hfe;
s_mem_contents[14'h1500] = 8'h68;
s_mem_contents[14'h1501] = 8'h49;
s_mem_contents[14'h1502] = 8'h30;
s_mem_contents[14'h1503] = 8'hcd;
s_mem_contents[14'h1504] = 8'h1d;
s_mem_contents[14'h1505] = 8'h02;
s_mem_contents[14'h1506] = 8'hd0;
s_mem_contents[14'h1507] = 8'hfe;
s_mem_contents[14'h1508] = 8'ha9;
s_mem_contents[14'h1509] = 8'h00;
s_mem_contents[14'h150a] = 8'h48;
s_mem_contents[14'h150b] = 8'h28;
s_mem_contents[14'h150c] = 8'ha0;
s_mem_contents[14'h150d] = 8'h41;
s_mem_contents[14'h150e] = 8'h08;
s_mem_contents[14'h150f] = 8'hcc;
s_mem_contents[14'h1510] = 8'h19;
s_mem_contents[14'h1511] = 8'h02;
s_mem_contents[14'h1512] = 8'hd0;
s_mem_contents[14'h1513] = 8'hfe;
s_mem_contents[14'h1514] = 8'h68;
s_mem_contents[14'h1515] = 8'h49;
s_mem_contents[14'h1516] = 8'h30;
s_mem_contents[14'h1517] = 8'hcd;
s_mem_contents[14'h1518] = 8'h1e;
s_mem_contents[14'h1519] = 8'h02;
s_mem_contents[14'h151a] = 8'hd0;
s_mem_contents[14'h151b] = 8'hfe;
s_mem_contents[14'h151c] = 8'ha9;
s_mem_contents[14'h151d] = 8'h00;
s_mem_contents[14'h151e] = 8'h48;
s_mem_contents[14'h151f] = 8'h28;
s_mem_contents[14'h1520] = 8'ha0;
s_mem_contents[14'h1521] = 8'h00;
s_mem_contents[14'h1522] = 8'h08;
s_mem_contents[14'h1523] = 8'hcc;
s_mem_contents[14'h1524] = 8'h1a;
s_mem_contents[14'h1525] = 8'h02;
s_mem_contents[14'h1526] = 8'hd0;
s_mem_contents[14'h1527] = 8'hfe;
s_mem_contents[14'h1528] = 8'h68;
s_mem_contents[14'h1529] = 8'h49;
s_mem_contents[14'h152a] = 8'h30;
s_mem_contents[14'h152b] = 8'hcd;
s_mem_contents[14'h152c] = 8'h1f;
s_mem_contents[14'h152d] = 8'h02;
s_mem_contents[14'h152e] = 8'hd0;
s_mem_contents[14'h152f] = 8'hfe;
s_mem_contents[14'h1530] = 8'ha9;
s_mem_contents[14'h1531] = 8'hff;
s_mem_contents[14'h1532] = 8'h48;
s_mem_contents[14'h1533] = 8'h28;
s_mem_contents[14'h1534] = 8'ha0;
s_mem_contents[14'h1535] = 8'hc3;
s_mem_contents[14'h1536] = 8'h08;
s_mem_contents[14'h1537] = 8'hcc;
s_mem_contents[14'h1538] = 8'h17;
s_mem_contents[14'h1539] = 8'h02;
s_mem_contents[14'h153a] = 8'hd0;
s_mem_contents[14'h153b] = 8'hfe;
s_mem_contents[14'h153c] = 8'h68;
s_mem_contents[14'h153d] = 8'h49;
s_mem_contents[14'h153e] = 8'h7d;
s_mem_contents[14'h153f] = 8'hcd;
s_mem_contents[14'h1540] = 8'h1c;
s_mem_contents[14'h1541] = 8'h02;
s_mem_contents[14'h1542] = 8'hd0;
s_mem_contents[14'h1543] = 8'hfe;
s_mem_contents[14'h1544] = 8'ha9;
s_mem_contents[14'h1545] = 8'hff;
s_mem_contents[14'h1546] = 8'h48;
s_mem_contents[14'h1547] = 8'h28;
s_mem_contents[14'h1548] = 8'ha0;
s_mem_contents[14'h1549] = 8'h82;
s_mem_contents[14'h154a] = 8'h08;
s_mem_contents[14'h154b] = 8'hcc;
s_mem_contents[14'h154c] = 8'h18;
s_mem_contents[14'h154d] = 8'h02;
s_mem_contents[14'h154e] = 8'hd0;
s_mem_contents[14'h154f] = 8'hfe;
s_mem_contents[14'h1550] = 8'h68;
s_mem_contents[14'h1551] = 8'h49;
s_mem_contents[14'h1552] = 8'h7d;
s_mem_contents[14'h1553] = 8'hcd;
s_mem_contents[14'h1554] = 8'h1d;
s_mem_contents[14'h1555] = 8'h02;
s_mem_contents[14'h1556] = 8'hd0;
s_mem_contents[14'h1557] = 8'hfe;
s_mem_contents[14'h1558] = 8'ha9;
s_mem_contents[14'h1559] = 8'hff;
s_mem_contents[14'h155a] = 8'h48;
s_mem_contents[14'h155b] = 8'h28;
s_mem_contents[14'h155c] = 8'ha0;
s_mem_contents[14'h155d] = 8'h41;
s_mem_contents[14'h155e] = 8'h08;
s_mem_contents[14'h155f] = 8'hcc;
s_mem_contents[14'h1560] = 8'h19;
s_mem_contents[14'h1561] = 8'h02;
s_mem_contents[14'h1562] = 8'hd0;
s_mem_contents[14'h1563] = 8'hfe;
s_mem_contents[14'h1564] = 8'h68;
s_mem_contents[14'h1565] = 8'h49;
s_mem_contents[14'h1566] = 8'h7d;
s_mem_contents[14'h1567] = 8'hcd;
s_mem_contents[14'h1568] = 8'h1e;
s_mem_contents[14'h1569] = 8'h02;
s_mem_contents[14'h156a] = 8'hd0;
s_mem_contents[14'h156b] = 8'hfe;
s_mem_contents[14'h156c] = 8'ha9;
s_mem_contents[14'h156d] = 8'hff;
s_mem_contents[14'h156e] = 8'h48;
s_mem_contents[14'h156f] = 8'h28;
s_mem_contents[14'h1570] = 8'ha0;
s_mem_contents[14'h1571] = 8'h00;
s_mem_contents[14'h1572] = 8'h08;
s_mem_contents[14'h1573] = 8'hcc;
s_mem_contents[14'h1574] = 8'h1a;
s_mem_contents[14'h1575] = 8'h02;
s_mem_contents[14'h1576] = 8'hd0;
s_mem_contents[14'h1577] = 8'hfe;
s_mem_contents[14'h1578] = 8'h68;
s_mem_contents[14'h1579] = 8'h49;
s_mem_contents[14'h157a] = 8'h7d;
s_mem_contents[14'h157b] = 8'hcd;
s_mem_contents[14'h157c] = 8'h1f;
s_mem_contents[14'h157d] = 8'h02;
s_mem_contents[14'h157e] = 8'hd0;
s_mem_contents[14'h157f] = 8'hfe;
s_mem_contents[14'h1580] = 8'ha0;
s_mem_contents[14'h1581] = 8'h00;
s_mem_contents[14'h1582] = 8'ha5;
s_mem_contents[14'h1583] = 8'h02;
s_mem_contents[14'h1584] = 8'h49;
s_mem_contents[14'h1585] = 8'hc3;
s_mem_contents[14'h1586] = 8'hc5;
s_mem_contents[14'h1587] = 8'h09;
s_mem_contents[14'h1588] = 8'hd0;
s_mem_contents[14'h1589] = 8'hfe;
s_mem_contents[14'h158a] = 8'h84;
s_mem_contents[14'h158b] = 8'h02;
s_mem_contents[14'h158c] = 8'had;
s_mem_contents[14'h158d] = 8'h03;
s_mem_contents[14'h158e] = 8'h02;
s_mem_contents[14'h158f] = 8'h49;
s_mem_contents[14'h1590] = 8'hc3;
s_mem_contents[14'h1591] = 8'hcd;
s_mem_contents[14'h1592] = 8'h17;
s_mem_contents[14'h1593] = 8'h02;
s_mem_contents[14'h1594] = 8'hd0;
s_mem_contents[14'h1595] = 8'hfe;
s_mem_contents[14'h1596] = 8'h8c;
s_mem_contents[14'h1597] = 8'h03;
s_mem_contents[14'h1598] = 8'h02;
s_mem_contents[14'h1599] = 8'ha5;
s_mem_contents[14'h159a] = 8'h03;
s_mem_contents[14'h159b] = 8'h49;
s_mem_contents[14'h159c] = 8'hc3;
s_mem_contents[14'h159d] = 8'hc5;
s_mem_contents[14'h159e] = 8'h0a;
s_mem_contents[14'h159f] = 8'hd0;
s_mem_contents[14'h15a0] = 8'hfe;
s_mem_contents[14'h15a1] = 8'h84;
s_mem_contents[14'h15a2] = 8'h03;
s_mem_contents[14'h15a3] = 8'had;
s_mem_contents[14'h15a4] = 8'h04;
s_mem_contents[14'h15a5] = 8'h02;
s_mem_contents[14'h15a6] = 8'h49;
s_mem_contents[14'h15a7] = 8'hc3;
s_mem_contents[14'h15a8] = 8'hcd;
s_mem_contents[14'h15a9] = 8'h18;
s_mem_contents[14'h15aa] = 8'h02;
s_mem_contents[14'h15ab] = 8'hd0;
s_mem_contents[14'h15ac] = 8'hfe;
s_mem_contents[14'h15ad] = 8'h8c;
s_mem_contents[14'h15ae] = 8'h04;
s_mem_contents[14'h15af] = 8'h02;
s_mem_contents[14'h15b0] = 8'ha5;
s_mem_contents[14'h15b1] = 8'h04;
s_mem_contents[14'h15b2] = 8'h49;
s_mem_contents[14'h15b3] = 8'hc3;
s_mem_contents[14'h15b4] = 8'hc5;
s_mem_contents[14'h15b5] = 8'h0b;
s_mem_contents[14'h15b6] = 8'hd0;
s_mem_contents[14'h15b7] = 8'hfe;
s_mem_contents[14'h15b8] = 8'h84;
s_mem_contents[14'h15b9] = 8'h04;
s_mem_contents[14'h15ba] = 8'had;
s_mem_contents[14'h15bb] = 8'h05;
s_mem_contents[14'h15bc] = 8'h02;
s_mem_contents[14'h15bd] = 8'h49;
s_mem_contents[14'h15be] = 8'hc3;
s_mem_contents[14'h15bf] = 8'hcd;
s_mem_contents[14'h15c0] = 8'h19;
s_mem_contents[14'h15c1] = 8'h02;
s_mem_contents[14'h15c2] = 8'hd0;
s_mem_contents[14'h15c3] = 8'hfe;
s_mem_contents[14'h15c4] = 8'h8c;
s_mem_contents[14'h15c5] = 8'h05;
s_mem_contents[14'h15c6] = 8'h02;
s_mem_contents[14'h15c7] = 8'ha5;
s_mem_contents[14'h15c8] = 8'h05;
s_mem_contents[14'h15c9] = 8'h49;
s_mem_contents[14'h15ca] = 8'hc3;
s_mem_contents[14'h15cb] = 8'hc5;
s_mem_contents[14'h15cc] = 8'h0c;
s_mem_contents[14'h15cd] = 8'hd0;
s_mem_contents[14'h15ce] = 8'hfe;
s_mem_contents[14'h15cf] = 8'h84;
s_mem_contents[14'h15d0] = 8'h05;
s_mem_contents[14'h15d1] = 8'had;
s_mem_contents[14'h15d2] = 8'h06;
s_mem_contents[14'h15d3] = 8'h02;
s_mem_contents[14'h15d4] = 8'h49;
s_mem_contents[14'h15d5] = 8'hc3;
s_mem_contents[14'h15d6] = 8'hcd;
s_mem_contents[14'h15d7] = 8'h1a;
s_mem_contents[14'h15d8] = 8'h02;
s_mem_contents[14'h15d9] = 8'hd0;
s_mem_contents[14'h15da] = 8'hfe;
s_mem_contents[14'h15db] = 8'h8c;
s_mem_contents[14'h15dc] = 8'h06;
s_mem_contents[14'h15dd] = 8'h02;
s_mem_contents[14'h15de] = 8'had;
s_mem_contents[14'h15df] = 8'h00;
s_mem_contents[14'h15e0] = 8'h02;
s_mem_contents[14'h15e1] = 8'hc9;
s_mem_contents[14'h15e2] = 8'h14;
s_mem_contents[14'h15e3] = 8'hd0;
s_mem_contents[14'h15e4] = 8'hfe;
s_mem_contents[14'h15e5] = 8'ha9;
s_mem_contents[14'h15e6] = 8'h15;
s_mem_contents[14'h15e7] = 8'h8d;
s_mem_contents[14'h15e8] = 8'h00;
s_mem_contents[14'h15e9] = 8'h02;
s_mem_contents[14'h15ea] = 8'ha2;
s_mem_contents[14'h15eb] = 8'h03;
s_mem_contents[14'h15ec] = 8'ha9;
s_mem_contents[14'h15ed] = 8'h00;
s_mem_contents[14'h15ee] = 8'h48;
s_mem_contents[14'h15ef] = 8'h28;
s_mem_contents[14'h15f0] = 8'hb5;
s_mem_contents[14'h15f1] = 8'h09;
s_mem_contents[14'h15f2] = 8'h08;
s_mem_contents[14'h15f3] = 8'h49;
s_mem_contents[14'h15f4] = 8'hc3;
s_mem_contents[14'h15f5] = 8'h28;
s_mem_contents[14'h15f6] = 8'h9d;
s_mem_contents[14'h15f7] = 8'h03;
s_mem_contents[14'h15f8] = 8'h02;
s_mem_contents[14'h15f9] = 8'h08;
s_mem_contents[14'h15fa] = 8'h49;
s_mem_contents[14'h15fb] = 8'hc3;
s_mem_contents[14'h15fc] = 8'hdd;
s_mem_contents[14'h15fd] = 8'h17;
s_mem_contents[14'h15fe] = 8'h02;
s_mem_contents[14'h15ff] = 8'hd0;
s_mem_contents[14'h1600] = 8'hfe;
s_mem_contents[14'h1601] = 8'h68;
s_mem_contents[14'h1602] = 8'h49;
s_mem_contents[14'h1603] = 8'h30;
s_mem_contents[14'h1604] = 8'hdd;
s_mem_contents[14'h1605] = 8'h1c;
s_mem_contents[14'h1606] = 8'h02;
s_mem_contents[14'h1607] = 8'hd0;
s_mem_contents[14'h1608] = 8'hfe;
s_mem_contents[14'h1609] = 8'hca;
s_mem_contents[14'h160a] = 8'h10;
s_mem_contents[14'h160b] = 8'he0;
s_mem_contents[14'h160c] = 8'ha2;
s_mem_contents[14'h160d] = 8'h03;
s_mem_contents[14'h160e] = 8'ha9;
s_mem_contents[14'h160f] = 8'hff;
s_mem_contents[14'h1610] = 8'h48;
s_mem_contents[14'h1611] = 8'h28;
s_mem_contents[14'h1612] = 8'hb5;
s_mem_contents[14'h1613] = 8'h09;
s_mem_contents[14'h1614] = 8'h08;
s_mem_contents[14'h1615] = 8'h49;
s_mem_contents[14'h1616] = 8'hc3;
s_mem_contents[14'h1617] = 8'h28;
s_mem_contents[14'h1618] = 8'h9d;
s_mem_contents[14'h1619] = 8'h03;
s_mem_contents[14'h161a] = 8'h02;
s_mem_contents[14'h161b] = 8'h08;
s_mem_contents[14'h161c] = 8'h49;
s_mem_contents[14'h161d] = 8'hc3;
s_mem_contents[14'h161e] = 8'hdd;
s_mem_contents[14'h161f] = 8'h17;
s_mem_contents[14'h1620] = 8'h02;
s_mem_contents[14'h1621] = 8'hd0;
s_mem_contents[14'h1622] = 8'hfe;
s_mem_contents[14'h1623] = 8'h68;
s_mem_contents[14'h1624] = 8'h49;
s_mem_contents[14'h1625] = 8'h7d;
s_mem_contents[14'h1626] = 8'hdd;
s_mem_contents[14'h1627] = 8'h1c;
s_mem_contents[14'h1628] = 8'h02;
s_mem_contents[14'h1629] = 8'hd0;
s_mem_contents[14'h162a] = 8'hfe;
s_mem_contents[14'h162b] = 8'hca;
s_mem_contents[14'h162c] = 8'h10;
s_mem_contents[14'h162d] = 8'he0;
s_mem_contents[14'h162e] = 8'ha2;
s_mem_contents[14'h162f] = 8'h03;
s_mem_contents[14'h1630] = 8'ha9;
s_mem_contents[14'h1631] = 8'h00;
s_mem_contents[14'h1632] = 8'h48;
s_mem_contents[14'h1633] = 8'h28;
s_mem_contents[14'h1634] = 8'hbd;
s_mem_contents[14'h1635] = 8'h17;
s_mem_contents[14'h1636] = 8'h02;
s_mem_contents[14'h1637] = 8'h08;
s_mem_contents[14'h1638] = 8'h49;
s_mem_contents[14'h1639] = 8'hc3;
s_mem_contents[14'h163a] = 8'h28;
s_mem_contents[14'h163b] = 8'h95;
s_mem_contents[14'h163c] = 8'h02;
s_mem_contents[14'h163d] = 8'h08;
s_mem_contents[14'h163e] = 8'h49;
s_mem_contents[14'h163f] = 8'hc3;
s_mem_contents[14'h1640] = 8'hd5;
s_mem_contents[14'h1641] = 8'h09;
s_mem_contents[14'h1642] = 8'hd0;
s_mem_contents[14'h1643] = 8'hfe;
s_mem_contents[14'h1644] = 8'h68;
s_mem_contents[14'h1645] = 8'h49;
s_mem_contents[14'h1646] = 8'h30;
s_mem_contents[14'h1647] = 8'hdd;
s_mem_contents[14'h1648] = 8'h1c;
s_mem_contents[14'h1649] = 8'h02;
s_mem_contents[14'h164a] = 8'hd0;
s_mem_contents[14'h164b] = 8'hfe;
s_mem_contents[14'h164c] = 8'hca;
s_mem_contents[14'h164d] = 8'h10;
s_mem_contents[14'h164e] = 8'he1;
s_mem_contents[14'h164f] = 8'ha2;
s_mem_contents[14'h1650] = 8'h03;
s_mem_contents[14'h1651] = 8'ha9;
s_mem_contents[14'h1652] = 8'hff;
s_mem_contents[14'h1653] = 8'h48;
s_mem_contents[14'h1654] = 8'h28;
s_mem_contents[14'h1655] = 8'hbd;
s_mem_contents[14'h1656] = 8'h17;
s_mem_contents[14'h1657] = 8'h02;
s_mem_contents[14'h1658] = 8'h08;
s_mem_contents[14'h1659] = 8'h49;
s_mem_contents[14'h165a] = 8'hc3;
s_mem_contents[14'h165b] = 8'h28;
s_mem_contents[14'h165c] = 8'h95;
s_mem_contents[14'h165d] = 8'h02;
s_mem_contents[14'h165e] = 8'h08;
s_mem_contents[14'h165f] = 8'h49;
s_mem_contents[14'h1660] = 8'hc3;
s_mem_contents[14'h1661] = 8'hd5;
s_mem_contents[14'h1662] = 8'h09;
s_mem_contents[14'h1663] = 8'hd0;
s_mem_contents[14'h1664] = 8'hfe;
s_mem_contents[14'h1665] = 8'h68;
s_mem_contents[14'h1666] = 8'h49;
s_mem_contents[14'h1667] = 8'h7d;
s_mem_contents[14'h1668] = 8'hdd;
s_mem_contents[14'h1669] = 8'h1c;
s_mem_contents[14'h166a] = 8'h02;
s_mem_contents[14'h166b] = 8'hd0;
s_mem_contents[14'h166c] = 8'hfe;
s_mem_contents[14'h166d] = 8'hca;
s_mem_contents[14'h166e] = 8'h10;
s_mem_contents[14'h166f] = 8'he1;
s_mem_contents[14'h1670] = 8'ha2;
s_mem_contents[14'h1671] = 8'h03;
s_mem_contents[14'h1672] = 8'ha0;
s_mem_contents[14'h1673] = 8'h00;
s_mem_contents[14'h1674] = 8'hb5;
s_mem_contents[14'h1675] = 8'h02;
s_mem_contents[14'h1676] = 8'h49;
s_mem_contents[14'h1677] = 8'hc3;
s_mem_contents[14'h1678] = 8'hd5;
s_mem_contents[14'h1679] = 8'h09;
s_mem_contents[14'h167a] = 8'hd0;
s_mem_contents[14'h167b] = 8'hfe;
s_mem_contents[14'h167c] = 8'h94;
s_mem_contents[14'h167d] = 8'h02;
s_mem_contents[14'h167e] = 8'hbd;
s_mem_contents[14'h167f] = 8'h03;
s_mem_contents[14'h1680] = 8'h02;
s_mem_contents[14'h1681] = 8'h49;
s_mem_contents[14'h1682] = 8'hc3;
s_mem_contents[14'h1683] = 8'hdd;
s_mem_contents[14'h1684] = 8'h17;
s_mem_contents[14'h1685] = 8'h02;
s_mem_contents[14'h1686] = 8'hd0;
s_mem_contents[14'h1687] = 8'hfe;
s_mem_contents[14'h1688] = 8'h8a;
s_mem_contents[14'h1689] = 8'h9d;
s_mem_contents[14'h168a] = 8'h03;
s_mem_contents[14'h168b] = 8'h02;
s_mem_contents[14'h168c] = 8'hca;
s_mem_contents[14'h168d] = 8'h10;
s_mem_contents[14'h168e] = 8'he5;
s_mem_contents[14'h168f] = 8'had;
s_mem_contents[14'h1690] = 8'h00;
s_mem_contents[14'h1691] = 8'h02;
s_mem_contents[14'h1692] = 8'hc9;
s_mem_contents[14'h1693] = 8'h15;
s_mem_contents[14'h1694] = 8'hd0;
s_mem_contents[14'h1695] = 8'hfe;
s_mem_contents[14'h1696] = 8'ha9;
s_mem_contents[14'h1697] = 8'h16;
s_mem_contents[14'h1698] = 8'h8d;
s_mem_contents[14'h1699] = 8'h00;
s_mem_contents[14'h169a] = 8'h02;
s_mem_contents[14'h169b] = 8'ha0;
s_mem_contents[14'h169c] = 8'h03;
s_mem_contents[14'h169d] = 8'ha9;
s_mem_contents[14'h169e] = 8'h00;
s_mem_contents[14'h169f] = 8'h48;
s_mem_contents[14'h16a0] = 8'h28;
s_mem_contents[14'h16a1] = 8'hb1;
s_mem_contents[14'h16a2] = 8'h1a;
s_mem_contents[14'h16a3] = 8'h08;
s_mem_contents[14'h16a4] = 8'h49;
s_mem_contents[14'h16a5] = 8'hc3;
s_mem_contents[14'h16a6] = 8'h28;
s_mem_contents[14'h16a7] = 8'h99;
s_mem_contents[14'h16a8] = 8'h03;
s_mem_contents[14'h16a9] = 8'h02;
s_mem_contents[14'h16aa] = 8'h08;
s_mem_contents[14'h16ab] = 8'h49;
s_mem_contents[14'h16ac] = 8'hc3;
s_mem_contents[14'h16ad] = 8'hd9;
s_mem_contents[14'h16ae] = 8'h17;
s_mem_contents[14'h16af] = 8'h02;
s_mem_contents[14'h16b0] = 8'hd0;
s_mem_contents[14'h16b1] = 8'hfe;
s_mem_contents[14'h16b2] = 8'h68;
s_mem_contents[14'h16b3] = 8'h49;
s_mem_contents[14'h16b4] = 8'h30;
s_mem_contents[14'h16b5] = 8'hd9;
s_mem_contents[14'h16b6] = 8'h1c;
s_mem_contents[14'h16b7] = 8'h02;
s_mem_contents[14'h16b8] = 8'hd0;
s_mem_contents[14'h16b9] = 8'hfe;
s_mem_contents[14'h16ba] = 8'h88;
s_mem_contents[14'h16bb] = 8'h10;
s_mem_contents[14'h16bc] = 8'he0;
s_mem_contents[14'h16bd] = 8'ha0;
s_mem_contents[14'h16be] = 8'h03;
s_mem_contents[14'h16bf] = 8'ha9;
s_mem_contents[14'h16c0] = 8'hff;
s_mem_contents[14'h16c1] = 8'h48;
s_mem_contents[14'h16c2] = 8'h28;
s_mem_contents[14'h16c3] = 8'hb1;
s_mem_contents[14'h16c4] = 8'h1a;
s_mem_contents[14'h16c5] = 8'h08;
s_mem_contents[14'h16c6] = 8'h49;
s_mem_contents[14'h16c7] = 8'hc3;
s_mem_contents[14'h16c8] = 8'h28;
s_mem_contents[14'h16c9] = 8'h99;
s_mem_contents[14'h16ca] = 8'h03;
s_mem_contents[14'h16cb] = 8'h02;
s_mem_contents[14'h16cc] = 8'h08;
s_mem_contents[14'h16cd] = 8'h49;
s_mem_contents[14'h16ce] = 8'hc3;
s_mem_contents[14'h16cf] = 8'hd9;
s_mem_contents[14'h16d0] = 8'h17;
s_mem_contents[14'h16d1] = 8'h02;
s_mem_contents[14'h16d2] = 8'hd0;
s_mem_contents[14'h16d3] = 8'hfe;
s_mem_contents[14'h16d4] = 8'h68;
s_mem_contents[14'h16d5] = 8'h49;
s_mem_contents[14'h16d6] = 8'h7d;
s_mem_contents[14'h16d7] = 8'hd9;
s_mem_contents[14'h16d8] = 8'h1c;
s_mem_contents[14'h16d9] = 8'h02;
s_mem_contents[14'h16da] = 8'hd0;
s_mem_contents[14'h16db] = 8'hfe;
s_mem_contents[14'h16dc] = 8'h88;
s_mem_contents[14'h16dd] = 8'h10;
s_mem_contents[14'h16de] = 8'he0;
s_mem_contents[14'h16df] = 8'ha0;
s_mem_contents[14'h16e0] = 8'h03;
s_mem_contents[14'h16e1] = 8'ha2;
s_mem_contents[14'h16e2] = 8'h00;
s_mem_contents[14'h16e3] = 8'hb9;
s_mem_contents[14'h16e4] = 8'h03;
s_mem_contents[14'h16e5] = 8'h02;
s_mem_contents[14'h16e6] = 8'h49;
s_mem_contents[14'h16e7] = 8'hc3;
s_mem_contents[14'h16e8] = 8'hd9;
s_mem_contents[14'h16e9] = 8'h17;
s_mem_contents[14'h16ea] = 8'h02;
s_mem_contents[14'h16eb] = 8'hd0;
s_mem_contents[14'h16ec] = 8'hfe;
s_mem_contents[14'h16ed] = 8'h8a;
s_mem_contents[14'h16ee] = 8'h99;
s_mem_contents[14'h16ef] = 8'h03;
s_mem_contents[14'h16f0] = 8'h02;
s_mem_contents[14'h16f1] = 8'h88;
s_mem_contents[14'h16f2] = 8'h10;
s_mem_contents[14'h16f3] = 8'hef;
s_mem_contents[14'h16f4] = 8'ha0;
s_mem_contents[14'h16f5] = 8'h03;
s_mem_contents[14'h16f6] = 8'ha9;
s_mem_contents[14'h16f7] = 8'h00;
s_mem_contents[14'h16f8] = 8'h48;
s_mem_contents[14'h16f9] = 8'h28;
s_mem_contents[14'h16fa] = 8'hb9;
s_mem_contents[14'h16fb] = 8'h17;
s_mem_contents[14'h16fc] = 8'h02;
s_mem_contents[14'h16fd] = 8'h08;
s_mem_contents[14'h16fe] = 8'h49;
s_mem_contents[14'h16ff] = 8'hc3;
s_mem_contents[14'h1700] = 8'h28;
s_mem_contents[14'h1701] = 8'h91;
s_mem_contents[14'h1702] = 8'h26;
s_mem_contents[14'h1703] = 8'h08;
s_mem_contents[14'h1704] = 8'h49;
s_mem_contents[14'h1705] = 8'hc3;
s_mem_contents[14'h1706] = 8'hd1;
s_mem_contents[14'h1707] = 8'h1a;
s_mem_contents[14'h1708] = 8'hd0;
s_mem_contents[14'h1709] = 8'hfe;
s_mem_contents[14'h170a] = 8'h68;
s_mem_contents[14'h170b] = 8'h49;
s_mem_contents[14'h170c] = 8'h30;
s_mem_contents[14'h170d] = 8'hd9;
s_mem_contents[14'h170e] = 8'h1c;
s_mem_contents[14'h170f] = 8'h02;
s_mem_contents[14'h1710] = 8'hd0;
s_mem_contents[14'h1711] = 8'hfe;
s_mem_contents[14'h1712] = 8'h88;
s_mem_contents[14'h1713] = 8'h10;
s_mem_contents[14'h1714] = 8'he1;
s_mem_contents[14'h1715] = 8'ha0;
s_mem_contents[14'h1716] = 8'h03;
s_mem_contents[14'h1717] = 8'ha9;
s_mem_contents[14'h1718] = 8'hff;
s_mem_contents[14'h1719] = 8'h48;
s_mem_contents[14'h171a] = 8'h28;
s_mem_contents[14'h171b] = 8'hb9;
s_mem_contents[14'h171c] = 8'h17;
s_mem_contents[14'h171d] = 8'h02;
s_mem_contents[14'h171e] = 8'h08;
s_mem_contents[14'h171f] = 8'h49;
s_mem_contents[14'h1720] = 8'hc3;
s_mem_contents[14'h1721] = 8'h28;
s_mem_contents[14'h1722] = 8'h91;
s_mem_contents[14'h1723] = 8'h26;
s_mem_contents[14'h1724] = 8'h08;
s_mem_contents[14'h1725] = 8'h49;
s_mem_contents[14'h1726] = 8'hc3;
s_mem_contents[14'h1727] = 8'hd1;
s_mem_contents[14'h1728] = 8'h1a;
s_mem_contents[14'h1729] = 8'hd0;
s_mem_contents[14'h172a] = 8'hfe;
s_mem_contents[14'h172b] = 8'h68;
s_mem_contents[14'h172c] = 8'h49;
s_mem_contents[14'h172d] = 8'h7d;
s_mem_contents[14'h172e] = 8'hd9;
s_mem_contents[14'h172f] = 8'h1c;
s_mem_contents[14'h1730] = 8'h02;
s_mem_contents[14'h1731] = 8'hd0;
s_mem_contents[14'h1732] = 8'hfe;
s_mem_contents[14'h1733] = 8'h88;
s_mem_contents[14'h1734] = 8'h10;
s_mem_contents[14'h1735] = 8'he1;
s_mem_contents[14'h1736] = 8'ha0;
s_mem_contents[14'h1737] = 8'h03;
s_mem_contents[14'h1738] = 8'ha2;
s_mem_contents[14'h1739] = 8'h00;
s_mem_contents[14'h173a] = 8'hb9;
s_mem_contents[14'h173b] = 8'h03;
s_mem_contents[14'h173c] = 8'h02;
s_mem_contents[14'h173d] = 8'h49;
s_mem_contents[14'h173e] = 8'hc3;
s_mem_contents[14'h173f] = 8'hd9;
s_mem_contents[14'h1740] = 8'h17;
s_mem_contents[14'h1741] = 8'h02;
s_mem_contents[14'h1742] = 8'hd0;
s_mem_contents[14'h1743] = 8'hfe;
s_mem_contents[14'h1744] = 8'h8a;
s_mem_contents[14'h1745] = 8'h99;
s_mem_contents[14'h1746] = 8'h03;
s_mem_contents[14'h1747] = 8'h02;
s_mem_contents[14'h1748] = 8'h88;
s_mem_contents[14'h1749] = 8'h10;
s_mem_contents[14'h174a] = 8'hef;
s_mem_contents[14'h174b] = 8'ha2;
s_mem_contents[14'h174c] = 8'h06;
s_mem_contents[14'h174d] = 8'ha0;
s_mem_contents[14'h174e] = 8'h03;
s_mem_contents[14'h174f] = 8'ha9;
s_mem_contents[14'h1750] = 8'h00;
s_mem_contents[14'h1751] = 8'h48;
s_mem_contents[14'h1752] = 8'h28;
s_mem_contents[14'h1753] = 8'ha1;
s_mem_contents[14'h1754] = 8'h1a;
s_mem_contents[14'h1755] = 8'h08;
s_mem_contents[14'h1756] = 8'h49;
s_mem_contents[14'h1757] = 8'hc3;
s_mem_contents[14'h1758] = 8'h28;
s_mem_contents[14'h1759] = 8'h81;
s_mem_contents[14'h175a] = 8'h26;
s_mem_contents[14'h175b] = 8'h08;
s_mem_contents[14'h175c] = 8'h49;
s_mem_contents[14'h175d] = 8'hc3;
s_mem_contents[14'h175e] = 8'hd9;
s_mem_contents[14'h175f] = 8'h17;
s_mem_contents[14'h1760] = 8'h02;
s_mem_contents[14'h1761] = 8'hd0;
s_mem_contents[14'h1762] = 8'hfe;
s_mem_contents[14'h1763] = 8'h68;
s_mem_contents[14'h1764] = 8'h49;
s_mem_contents[14'h1765] = 8'h30;
s_mem_contents[14'h1766] = 8'hd9;
s_mem_contents[14'h1767] = 8'h1c;
s_mem_contents[14'h1768] = 8'h02;
s_mem_contents[14'h1769] = 8'hd0;
s_mem_contents[14'h176a] = 8'hfe;
s_mem_contents[14'h176b] = 8'hca;
s_mem_contents[14'h176c] = 8'hca;
s_mem_contents[14'h176d] = 8'h88;
s_mem_contents[14'h176e] = 8'h10;
s_mem_contents[14'h176f] = 8'hdf;
s_mem_contents[14'h1770] = 8'ha2;
s_mem_contents[14'h1771] = 8'h06;
s_mem_contents[14'h1772] = 8'ha0;
s_mem_contents[14'h1773] = 8'h03;
s_mem_contents[14'h1774] = 8'ha9;
s_mem_contents[14'h1775] = 8'hff;
s_mem_contents[14'h1776] = 8'h48;
s_mem_contents[14'h1777] = 8'h28;
s_mem_contents[14'h1778] = 8'ha1;
s_mem_contents[14'h1779] = 8'h1a;
s_mem_contents[14'h177a] = 8'h08;
s_mem_contents[14'h177b] = 8'h49;
s_mem_contents[14'h177c] = 8'hc3;
s_mem_contents[14'h177d] = 8'h28;
s_mem_contents[14'h177e] = 8'h81;
s_mem_contents[14'h177f] = 8'h26;
s_mem_contents[14'h1780] = 8'h08;
s_mem_contents[14'h1781] = 8'h49;
s_mem_contents[14'h1782] = 8'hc3;
s_mem_contents[14'h1783] = 8'hd9;
s_mem_contents[14'h1784] = 8'h17;
s_mem_contents[14'h1785] = 8'h02;
s_mem_contents[14'h1786] = 8'hd0;
s_mem_contents[14'h1787] = 8'hfe;
s_mem_contents[14'h1788] = 8'h68;
s_mem_contents[14'h1789] = 8'h49;
s_mem_contents[14'h178a] = 8'h7d;
s_mem_contents[14'h178b] = 8'hd9;
s_mem_contents[14'h178c] = 8'h1c;
s_mem_contents[14'h178d] = 8'h02;
s_mem_contents[14'h178e] = 8'hd0;
s_mem_contents[14'h178f] = 8'hfe;
s_mem_contents[14'h1790] = 8'hca;
s_mem_contents[14'h1791] = 8'hca;
s_mem_contents[14'h1792] = 8'h88;
s_mem_contents[14'h1793] = 8'h10;
s_mem_contents[14'h1794] = 8'hdf;
s_mem_contents[14'h1795] = 8'ha0;
s_mem_contents[14'h1796] = 8'h03;
s_mem_contents[14'h1797] = 8'ha2;
s_mem_contents[14'h1798] = 8'h00;
s_mem_contents[14'h1799] = 8'hb9;
s_mem_contents[14'h179a] = 8'h03;
s_mem_contents[14'h179b] = 8'h02;
s_mem_contents[14'h179c] = 8'h49;
s_mem_contents[14'h179d] = 8'hc3;
s_mem_contents[14'h179e] = 8'hd9;
s_mem_contents[14'h179f] = 8'h17;
s_mem_contents[14'h17a0] = 8'h02;
s_mem_contents[14'h17a1] = 8'hd0;
s_mem_contents[14'h17a2] = 8'hfe;
s_mem_contents[14'h17a3] = 8'h8a;
s_mem_contents[14'h17a4] = 8'h99;
s_mem_contents[14'h17a5] = 8'h03;
s_mem_contents[14'h17a6] = 8'h02;
s_mem_contents[14'h17a7] = 8'h88;
s_mem_contents[14'h17a8] = 8'h10;
s_mem_contents[14'h17a9] = 8'hef;
s_mem_contents[14'h17aa] = 8'had;
s_mem_contents[14'h17ab] = 8'h00;
s_mem_contents[14'h17ac] = 8'h02;
s_mem_contents[14'h17ad] = 8'hc9;
s_mem_contents[14'h17ae] = 8'h16;
s_mem_contents[14'h17af] = 8'hd0;
s_mem_contents[14'h17b0] = 8'hfe;
s_mem_contents[14'h17b1] = 8'ha9;
s_mem_contents[14'h17b2] = 8'h17;
s_mem_contents[14'h17b3] = 8'h8d;
s_mem_contents[14'h17b4] = 8'h00;
s_mem_contents[14'h17b5] = 8'h02;
s_mem_contents[14'h17b6] = 8'ha2;
s_mem_contents[14'h17b7] = 8'hfd;
s_mem_contents[14'h17b8] = 8'hb5;
s_mem_contents[14'h17b9] = 8'h0f;
s_mem_contents[14'h17ba] = 8'h9d;
s_mem_contents[14'h17bb] = 8'h09;
s_mem_contents[14'h17bc] = 8'h01;
s_mem_contents[14'h17bd] = 8'hca;
s_mem_contents[14'h17be] = 8'he0;
s_mem_contents[14'h17bf] = 8'hfa;
s_mem_contents[14'h17c0] = 8'hb0;
s_mem_contents[14'h17c1] = 8'hf6;
s_mem_contents[14'h17c2] = 8'ha2;
s_mem_contents[14'h17c3] = 8'hfd;
s_mem_contents[14'h17c4] = 8'hbd;
s_mem_contents[14'h17c5] = 8'h1d;
s_mem_contents[14'h17c6] = 8'h01;
s_mem_contents[14'h17c7] = 8'h95;
s_mem_contents[14'h17c8] = 8'h08;
s_mem_contents[14'h17c9] = 8'hca;
s_mem_contents[14'h17ca] = 8'he0;
s_mem_contents[14'h17cb] = 8'hfa;
s_mem_contents[14'h17cc] = 8'hb0;
s_mem_contents[14'h17cd] = 8'hf6;
s_mem_contents[14'h17ce] = 8'ha2;
s_mem_contents[14'h17cf] = 8'h03;
s_mem_contents[14'h17d0] = 8'ha0;
s_mem_contents[14'h17d1] = 8'h00;
s_mem_contents[14'h17d2] = 8'hb5;
s_mem_contents[14'h17d3] = 8'h02;
s_mem_contents[14'h17d4] = 8'hd5;
s_mem_contents[14'h17d5] = 8'h09;
s_mem_contents[14'h17d6] = 8'hd0;
s_mem_contents[14'h17d7] = 8'hfe;
s_mem_contents[14'h17d8] = 8'h94;
s_mem_contents[14'h17d9] = 8'h02;
s_mem_contents[14'h17da] = 8'hbd;
s_mem_contents[14'h17db] = 8'h03;
s_mem_contents[14'h17dc] = 8'h02;
s_mem_contents[14'h17dd] = 8'hdd;
s_mem_contents[14'h17de] = 8'h17;
s_mem_contents[14'h17df] = 8'h02;
s_mem_contents[14'h17e0] = 8'hd0;
s_mem_contents[14'h17e1] = 8'hfe;
s_mem_contents[14'h17e2] = 8'h8a;
s_mem_contents[14'h17e3] = 8'h9d;
s_mem_contents[14'h17e4] = 8'h03;
s_mem_contents[14'h17e5] = 8'h02;
s_mem_contents[14'h17e6] = 8'hca;
s_mem_contents[14'h17e7] = 8'h10;
s_mem_contents[14'h17e8] = 8'he9;
s_mem_contents[14'h17e9] = 8'ha0;
s_mem_contents[14'h17ea] = 8'hfb;
s_mem_contents[14'h17eb] = 8'ha2;
s_mem_contents[14'h17ec] = 8'hfe;
s_mem_contents[14'h17ed] = 8'ha1;
s_mem_contents[14'h17ee] = 8'h22;
s_mem_contents[14'h17ef] = 8'h99;
s_mem_contents[14'h17f0] = 8'h0b;
s_mem_contents[14'h17f1] = 8'h01;
s_mem_contents[14'h17f2] = 8'hca;
s_mem_contents[14'h17f3] = 8'hca;
s_mem_contents[14'h17f4] = 8'h88;
s_mem_contents[14'h17f5] = 8'hc0;
s_mem_contents[14'h17f6] = 8'hf8;
s_mem_contents[14'h17f7] = 8'hb0;
s_mem_contents[14'h17f8] = 8'hf4;
s_mem_contents[14'h17f9] = 8'ha0;
s_mem_contents[14'h17fa] = 8'h03;
s_mem_contents[14'h17fb] = 8'ha2;
s_mem_contents[14'h17fc] = 8'h00;
s_mem_contents[14'h17fd] = 8'hb9;
s_mem_contents[14'h17fe] = 8'h03;
s_mem_contents[14'h17ff] = 8'h02;
s_mem_contents[14'h1800] = 8'hd9;
s_mem_contents[14'h1801] = 8'h17;
s_mem_contents[14'h1802] = 8'h02;
s_mem_contents[14'h1803] = 8'hd0;
s_mem_contents[14'h1804] = 8'hfe;
s_mem_contents[14'h1805] = 8'h8a;
s_mem_contents[14'h1806] = 8'h99;
s_mem_contents[14'h1807] = 8'h03;
s_mem_contents[14'h1808] = 8'h02;
s_mem_contents[14'h1809] = 8'h88;
s_mem_contents[14'h180a] = 8'h10;
s_mem_contents[14'h180b] = 8'hf1;
s_mem_contents[14'h180c] = 8'ha0;
s_mem_contents[14'h180d] = 8'hfb;
s_mem_contents[14'h180e] = 8'hb9;
s_mem_contents[14'h180f] = 8'h1f;
s_mem_contents[14'h1810] = 8'h01;
s_mem_contents[14'h1811] = 8'h91;
s_mem_contents[14'h1812] = 8'h2e;
s_mem_contents[14'h1813] = 8'h88;
s_mem_contents[14'h1814] = 8'hc0;
s_mem_contents[14'h1815] = 8'hf8;
s_mem_contents[14'h1816] = 8'hb0;
s_mem_contents[14'h1817] = 8'hf6;
s_mem_contents[14'h1818] = 8'ha0;
s_mem_contents[14'h1819] = 8'h03;
s_mem_contents[14'h181a] = 8'ha2;
s_mem_contents[14'h181b] = 8'h00;
s_mem_contents[14'h181c] = 8'hb9;
s_mem_contents[14'h181d] = 8'h03;
s_mem_contents[14'h181e] = 8'h02;
s_mem_contents[14'h181f] = 8'hd9;
s_mem_contents[14'h1820] = 8'h17;
s_mem_contents[14'h1821] = 8'h02;
s_mem_contents[14'h1822] = 8'hd0;
s_mem_contents[14'h1823] = 8'hfe;
s_mem_contents[14'h1824] = 8'h8a;
s_mem_contents[14'h1825] = 8'h99;
s_mem_contents[14'h1826] = 8'h03;
s_mem_contents[14'h1827] = 8'h02;
s_mem_contents[14'h1828] = 8'h88;
s_mem_contents[14'h1829] = 8'h10;
s_mem_contents[14'h182a] = 8'hf1;
s_mem_contents[14'h182b] = 8'ha0;
s_mem_contents[14'h182c] = 8'hfb;
s_mem_contents[14'h182d] = 8'ha2;
s_mem_contents[14'h182e] = 8'hfe;
s_mem_contents[14'h182f] = 8'hb1;
s_mem_contents[14'h1830] = 8'h24;
s_mem_contents[14'h1831] = 8'h81;
s_mem_contents[14'h1832] = 8'h2e;
s_mem_contents[14'h1833] = 8'hca;
s_mem_contents[14'h1834] = 8'hca;
s_mem_contents[14'h1835] = 8'h88;
s_mem_contents[14'h1836] = 8'hc0;
s_mem_contents[14'h1837] = 8'hf8;
s_mem_contents[14'h1838] = 8'hb0;
s_mem_contents[14'h1839] = 8'hf5;
s_mem_contents[14'h183a] = 8'ha0;
s_mem_contents[14'h183b] = 8'h03;
s_mem_contents[14'h183c] = 8'ha2;
s_mem_contents[14'h183d] = 8'h00;
s_mem_contents[14'h183e] = 8'hb9;
s_mem_contents[14'h183f] = 8'h03;
s_mem_contents[14'h1840] = 8'h02;
s_mem_contents[14'h1841] = 8'hd9;
s_mem_contents[14'h1842] = 8'h17;
s_mem_contents[14'h1843] = 8'h02;
s_mem_contents[14'h1844] = 8'hd0;
s_mem_contents[14'h1845] = 8'hfe;
s_mem_contents[14'h1846] = 8'h8a;
s_mem_contents[14'h1847] = 8'h99;
s_mem_contents[14'h1848] = 8'h03;
s_mem_contents[14'h1849] = 8'h02;
s_mem_contents[14'h184a] = 8'h88;
s_mem_contents[14'h184b] = 8'h10;
s_mem_contents[14'h184c] = 8'hf1;
s_mem_contents[14'h184d] = 8'had;
s_mem_contents[14'h184e] = 8'h00;
s_mem_contents[14'h184f] = 8'h02;
s_mem_contents[14'h1850] = 8'hc9;
s_mem_contents[14'h1851] = 8'h17;
s_mem_contents[14'h1852] = 8'hd0;
s_mem_contents[14'h1853] = 8'hfe;
s_mem_contents[14'h1854] = 8'ha9;
s_mem_contents[14'h1855] = 8'h18;
s_mem_contents[14'h1856] = 8'h8d;
s_mem_contents[14'h1857] = 8'h00;
s_mem_contents[14'h1858] = 8'h02;
s_mem_contents[14'h1859] = 8'ha9;
s_mem_contents[14'h185a] = 8'h00;
s_mem_contents[14'h185b] = 8'h48;
s_mem_contents[14'h185c] = 8'h28;
s_mem_contents[14'h185d] = 8'ha5;
s_mem_contents[14'h185e] = 8'h09;
s_mem_contents[14'h185f] = 8'h08;
s_mem_contents[14'h1860] = 8'h49;
s_mem_contents[14'h1861] = 8'hc3;
s_mem_contents[14'h1862] = 8'h28;
s_mem_contents[14'h1863] = 8'h8d;
s_mem_contents[14'h1864] = 8'h03;
s_mem_contents[14'h1865] = 8'h02;
s_mem_contents[14'h1866] = 8'h08;
s_mem_contents[14'h1867] = 8'h49;
s_mem_contents[14'h1868] = 8'hc3;
s_mem_contents[14'h1869] = 8'hc9;
s_mem_contents[14'h186a] = 8'hc3;
s_mem_contents[14'h186b] = 8'hd0;
s_mem_contents[14'h186c] = 8'hfe;
s_mem_contents[14'h186d] = 8'h68;
s_mem_contents[14'h186e] = 8'h49;
s_mem_contents[14'h186f] = 8'h30;
s_mem_contents[14'h1870] = 8'hcd;
s_mem_contents[14'h1871] = 8'h1c;
s_mem_contents[14'h1872] = 8'h02;
s_mem_contents[14'h1873] = 8'hd0;
s_mem_contents[14'h1874] = 8'hfe;
s_mem_contents[14'h1875] = 8'ha9;
s_mem_contents[14'h1876] = 8'h00;
s_mem_contents[14'h1877] = 8'h48;
s_mem_contents[14'h1878] = 8'h28;
s_mem_contents[14'h1879] = 8'ha5;
s_mem_contents[14'h187a] = 8'h0a;
s_mem_contents[14'h187b] = 8'h08;
s_mem_contents[14'h187c] = 8'h49;
s_mem_contents[14'h187d] = 8'hc3;
s_mem_contents[14'h187e] = 8'h28;
s_mem_contents[14'h187f] = 8'h8d;
s_mem_contents[14'h1880] = 8'h04;
s_mem_contents[14'h1881] = 8'h02;
s_mem_contents[14'h1882] = 8'h08;
s_mem_contents[14'h1883] = 8'h49;
s_mem_contents[14'h1884] = 8'hc3;
s_mem_contents[14'h1885] = 8'hc9;
s_mem_contents[14'h1886] = 8'h82;
s_mem_contents[14'h1887] = 8'hd0;
s_mem_contents[14'h1888] = 8'hfe;
s_mem_contents[14'h1889] = 8'h68;
s_mem_contents[14'h188a] = 8'h49;
s_mem_contents[14'h188b] = 8'h30;
s_mem_contents[14'h188c] = 8'hcd;
s_mem_contents[14'h188d] = 8'h1d;
s_mem_contents[14'h188e] = 8'h02;
s_mem_contents[14'h188f] = 8'hd0;
s_mem_contents[14'h1890] = 8'hfe;
s_mem_contents[14'h1891] = 8'ha9;
s_mem_contents[14'h1892] = 8'h00;
s_mem_contents[14'h1893] = 8'h48;
s_mem_contents[14'h1894] = 8'h28;
s_mem_contents[14'h1895] = 8'ha5;
s_mem_contents[14'h1896] = 8'h0b;
s_mem_contents[14'h1897] = 8'h08;
s_mem_contents[14'h1898] = 8'h49;
s_mem_contents[14'h1899] = 8'hc3;
s_mem_contents[14'h189a] = 8'h28;
s_mem_contents[14'h189b] = 8'h8d;
s_mem_contents[14'h189c] = 8'h05;
s_mem_contents[14'h189d] = 8'h02;
s_mem_contents[14'h189e] = 8'h08;
s_mem_contents[14'h189f] = 8'h49;
s_mem_contents[14'h18a0] = 8'hc3;
s_mem_contents[14'h18a1] = 8'hc9;
s_mem_contents[14'h18a2] = 8'h41;
s_mem_contents[14'h18a3] = 8'hd0;
s_mem_contents[14'h18a4] = 8'hfe;
s_mem_contents[14'h18a5] = 8'h68;
s_mem_contents[14'h18a6] = 8'h49;
s_mem_contents[14'h18a7] = 8'h30;
s_mem_contents[14'h18a8] = 8'hcd;
s_mem_contents[14'h18a9] = 8'h1e;
s_mem_contents[14'h18aa] = 8'h02;
s_mem_contents[14'h18ab] = 8'hd0;
s_mem_contents[14'h18ac] = 8'hfe;
s_mem_contents[14'h18ad] = 8'ha9;
s_mem_contents[14'h18ae] = 8'h00;
s_mem_contents[14'h18af] = 8'h48;
s_mem_contents[14'h18b0] = 8'h28;
s_mem_contents[14'h18b1] = 8'ha5;
s_mem_contents[14'h18b2] = 8'h0c;
s_mem_contents[14'h18b3] = 8'h08;
s_mem_contents[14'h18b4] = 8'h49;
s_mem_contents[14'h18b5] = 8'hc3;
s_mem_contents[14'h18b6] = 8'h28;
s_mem_contents[14'h18b7] = 8'h8d;
s_mem_contents[14'h18b8] = 8'h06;
s_mem_contents[14'h18b9] = 8'h02;
s_mem_contents[14'h18ba] = 8'h08;
s_mem_contents[14'h18bb] = 8'h49;
s_mem_contents[14'h18bc] = 8'hc3;
s_mem_contents[14'h18bd] = 8'hc9;
s_mem_contents[14'h18be] = 8'h00;
s_mem_contents[14'h18bf] = 8'hd0;
s_mem_contents[14'h18c0] = 8'hfe;
s_mem_contents[14'h18c1] = 8'h68;
s_mem_contents[14'h18c2] = 8'h49;
s_mem_contents[14'h18c3] = 8'h30;
s_mem_contents[14'h18c4] = 8'hcd;
s_mem_contents[14'h18c5] = 8'h1f;
s_mem_contents[14'h18c6] = 8'h02;
s_mem_contents[14'h18c7] = 8'hd0;
s_mem_contents[14'h18c8] = 8'hfe;
s_mem_contents[14'h18c9] = 8'ha9;
s_mem_contents[14'h18ca] = 8'hff;
s_mem_contents[14'h18cb] = 8'h48;
s_mem_contents[14'h18cc] = 8'h28;
s_mem_contents[14'h18cd] = 8'ha5;
s_mem_contents[14'h18ce] = 8'h09;
s_mem_contents[14'h18cf] = 8'h08;
s_mem_contents[14'h18d0] = 8'h49;
s_mem_contents[14'h18d1] = 8'hc3;
s_mem_contents[14'h18d2] = 8'h28;
s_mem_contents[14'h18d3] = 8'h8d;
s_mem_contents[14'h18d4] = 8'h03;
s_mem_contents[14'h18d5] = 8'h02;
s_mem_contents[14'h18d6] = 8'h08;
s_mem_contents[14'h18d7] = 8'h49;
s_mem_contents[14'h18d8] = 8'hc3;
s_mem_contents[14'h18d9] = 8'hc9;
s_mem_contents[14'h18da] = 8'hc3;
s_mem_contents[14'h18db] = 8'hd0;
s_mem_contents[14'h18dc] = 8'hfe;
s_mem_contents[14'h18dd] = 8'h68;
s_mem_contents[14'h18de] = 8'h49;
s_mem_contents[14'h18df] = 8'h7d;
s_mem_contents[14'h18e0] = 8'hcd;
s_mem_contents[14'h18e1] = 8'h1c;
s_mem_contents[14'h18e2] = 8'h02;
s_mem_contents[14'h18e3] = 8'hd0;
s_mem_contents[14'h18e4] = 8'hfe;
s_mem_contents[14'h18e5] = 8'ha9;
s_mem_contents[14'h18e6] = 8'hff;
s_mem_contents[14'h18e7] = 8'h48;
s_mem_contents[14'h18e8] = 8'h28;
s_mem_contents[14'h18e9] = 8'ha5;
s_mem_contents[14'h18ea] = 8'h0a;
s_mem_contents[14'h18eb] = 8'h08;
s_mem_contents[14'h18ec] = 8'h49;
s_mem_contents[14'h18ed] = 8'hc3;
s_mem_contents[14'h18ee] = 8'h28;
s_mem_contents[14'h18ef] = 8'h8d;
s_mem_contents[14'h18f0] = 8'h04;
s_mem_contents[14'h18f1] = 8'h02;
s_mem_contents[14'h18f2] = 8'h08;
s_mem_contents[14'h18f3] = 8'h49;
s_mem_contents[14'h18f4] = 8'hc3;
s_mem_contents[14'h18f5] = 8'hc9;
s_mem_contents[14'h18f6] = 8'h82;
s_mem_contents[14'h18f7] = 8'hd0;
s_mem_contents[14'h18f8] = 8'hfe;
s_mem_contents[14'h18f9] = 8'h68;
s_mem_contents[14'h18fa] = 8'h49;
s_mem_contents[14'h18fb] = 8'h7d;
s_mem_contents[14'h18fc] = 8'hcd;
s_mem_contents[14'h18fd] = 8'h1d;
s_mem_contents[14'h18fe] = 8'h02;
s_mem_contents[14'h18ff] = 8'hd0;
s_mem_contents[14'h1900] = 8'hfe;
s_mem_contents[14'h1901] = 8'ha9;
s_mem_contents[14'h1902] = 8'hff;
s_mem_contents[14'h1903] = 8'h48;
s_mem_contents[14'h1904] = 8'h28;
s_mem_contents[14'h1905] = 8'ha5;
s_mem_contents[14'h1906] = 8'h0b;
s_mem_contents[14'h1907] = 8'h08;
s_mem_contents[14'h1908] = 8'h49;
s_mem_contents[14'h1909] = 8'hc3;
s_mem_contents[14'h190a] = 8'h28;
s_mem_contents[14'h190b] = 8'h8d;
s_mem_contents[14'h190c] = 8'h05;
s_mem_contents[14'h190d] = 8'h02;
s_mem_contents[14'h190e] = 8'h08;
s_mem_contents[14'h190f] = 8'h49;
s_mem_contents[14'h1910] = 8'hc3;
s_mem_contents[14'h1911] = 8'hc9;
s_mem_contents[14'h1912] = 8'h41;
s_mem_contents[14'h1913] = 8'hd0;
s_mem_contents[14'h1914] = 8'hfe;
s_mem_contents[14'h1915] = 8'h68;
s_mem_contents[14'h1916] = 8'h49;
s_mem_contents[14'h1917] = 8'h7d;
s_mem_contents[14'h1918] = 8'hcd;
s_mem_contents[14'h1919] = 8'h1e;
s_mem_contents[14'h191a] = 8'h02;
s_mem_contents[14'h191b] = 8'hd0;
s_mem_contents[14'h191c] = 8'hfe;
s_mem_contents[14'h191d] = 8'ha9;
s_mem_contents[14'h191e] = 8'hff;
s_mem_contents[14'h191f] = 8'h48;
s_mem_contents[14'h1920] = 8'h28;
s_mem_contents[14'h1921] = 8'ha5;
s_mem_contents[14'h1922] = 8'h0c;
s_mem_contents[14'h1923] = 8'h08;
s_mem_contents[14'h1924] = 8'h49;
s_mem_contents[14'h1925] = 8'hc3;
s_mem_contents[14'h1926] = 8'h28;
s_mem_contents[14'h1927] = 8'h8d;
s_mem_contents[14'h1928] = 8'h06;
s_mem_contents[14'h1929] = 8'h02;
s_mem_contents[14'h192a] = 8'h08;
s_mem_contents[14'h192b] = 8'h49;
s_mem_contents[14'h192c] = 8'hc3;
s_mem_contents[14'h192d] = 8'hc9;
s_mem_contents[14'h192e] = 8'h00;
s_mem_contents[14'h192f] = 8'hd0;
s_mem_contents[14'h1930] = 8'hfe;
s_mem_contents[14'h1931] = 8'h68;
s_mem_contents[14'h1932] = 8'h49;
s_mem_contents[14'h1933] = 8'h7d;
s_mem_contents[14'h1934] = 8'hcd;
s_mem_contents[14'h1935] = 8'h1f;
s_mem_contents[14'h1936] = 8'h02;
s_mem_contents[14'h1937] = 8'hd0;
s_mem_contents[14'h1938] = 8'hfe;
s_mem_contents[14'h1939] = 8'ha9;
s_mem_contents[14'h193a] = 8'h00;
s_mem_contents[14'h193b] = 8'h48;
s_mem_contents[14'h193c] = 8'h28;
s_mem_contents[14'h193d] = 8'had;
s_mem_contents[14'h193e] = 8'h17;
s_mem_contents[14'h193f] = 8'h02;
s_mem_contents[14'h1940] = 8'h08;
s_mem_contents[14'h1941] = 8'h49;
s_mem_contents[14'h1942] = 8'hc3;
s_mem_contents[14'h1943] = 8'h28;
s_mem_contents[14'h1944] = 8'h85;
s_mem_contents[14'h1945] = 8'h02;
s_mem_contents[14'h1946] = 8'h08;
s_mem_contents[14'h1947] = 8'h49;
s_mem_contents[14'h1948] = 8'hc3;
s_mem_contents[14'h1949] = 8'hc5;
s_mem_contents[14'h194a] = 8'h09;
s_mem_contents[14'h194b] = 8'hd0;
s_mem_contents[14'h194c] = 8'hfe;
s_mem_contents[14'h194d] = 8'h68;
s_mem_contents[14'h194e] = 8'h49;
s_mem_contents[14'h194f] = 8'h30;
s_mem_contents[14'h1950] = 8'hcd;
s_mem_contents[14'h1951] = 8'h1c;
s_mem_contents[14'h1952] = 8'h02;
s_mem_contents[14'h1953] = 8'hd0;
s_mem_contents[14'h1954] = 8'hfe;
s_mem_contents[14'h1955] = 8'ha9;
s_mem_contents[14'h1956] = 8'h00;
s_mem_contents[14'h1957] = 8'h48;
s_mem_contents[14'h1958] = 8'h28;
s_mem_contents[14'h1959] = 8'had;
s_mem_contents[14'h195a] = 8'h18;
s_mem_contents[14'h195b] = 8'h02;
s_mem_contents[14'h195c] = 8'h08;
s_mem_contents[14'h195d] = 8'h49;
s_mem_contents[14'h195e] = 8'hc3;
s_mem_contents[14'h195f] = 8'h28;
s_mem_contents[14'h1960] = 8'h85;
s_mem_contents[14'h1961] = 8'h03;
s_mem_contents[14'h1962] = 8'h08;
s_mem_contents[14'h1963] = 8'h49;
s_mem_contents[14'h1964] = 8'hc3;
s_mem_contents[14'h1965] = 8'hc5;
s_mem_contents[14'h1966] = 8'h0a;
s_mem_contents[14'h1967] = 8'hd0;
s_mem_contents[14'h1968] = 8'hfe;
s_mem_contents[14'h1969] = 8'h68;
s_mem_contents[14'h196a] = 8'h49;
s_mem_contents[14'h196b] = 8'h30;
s_mem_contents[14'h196c] = 8'hcd;
s_mem_contents[14'h196d] = 8'h1d;
s_mem_contents[14'h196e] = 8'h02;
s_mem_contents[14'h196f] = 8'hd0;
s_mem_contents[14'h1970] = 8'hfe;
s_mem_contents[14'h1971] = 8'ha9;
s_mem_contents[14'h1972] = 8'h00;
s_mem_contents[14'h1973] = 8'h48;
s_mem_contents[14'h1974] = 8'h28;
s_mem_contents[14'h1975] = 8'had;
s_mem_contents[14'h1976] = 8'h19;
s_mem_contents[14'h1977] = 8'h02;
s_mem_contents[14'h1978] = 8'h08;
s_mem_contents[14'h1979] = 8'h49;
s_mem_contents[14'h197a] = 8'hc3;
s_mem_contents[14'h197b] = 8'h28;
s_mem_contents[14'h197c] = 8'h85;
s_mem_contents[14'h197d] = 8'h04;
s_mem_contents[14'h197e] = 8'h08;
s_mem_contents[14'h197f] = 8'h49;
s_mem_contents[14'h1980] = 8'hc3;
s_mem_contents[14'h1981] = 8'hc5;
s_mem_contents[14'h1982] = 8'h0b;
s_mem_contents[14'h1983] = 8'hd0;
s_mem_contents[14'h1984] = 8'hfe;
s_mem_contents[14'h1985] = 8'h68;
s_mem_contents[14'h1986] = 8'h49;
s_mem_contents[14'h1987] = 8'h30;
s_mem_contents[14'h1988] = 8'hcd;
s_mem_contents[14'h1989] = 8'h1e;
s_mem_contents[14'h198a] = 8'h02;
s_mem_contents[14'h198b] = 8'hd0;
s_mem_contents[14'h198c] = 8'hfe;
s_mem_contents[14'h198d] = 8'ha9;
s_mem_contents[14'h198e] = 8'h00;
s_mem_contents[14'h198f] = 8'h48;
s_mem_contents[14'h1990] = 8'h28;
s_mem_contents[14'h1991] = 8'had;
s_mem_contents[14'h1992] = 8'h1a;
s_mem_contents[14'h1993] = 8'h02;
s_mem_contents[14'h1994] = 8'h08;
s_mem_contents[14'h1995] = 8'h49;
s_mem_contents[14'h1996] = 8'hc3;
s_mem_contents[14'h1997] = 8'h28;
s_mem_contents[14'h1998] = 8'h85;
s_mem_contents[14'h1999] = 8'h05;
s_mem_contents[14'h199a] = 8'h08;
s_mem_contents[14'h199b] = 8'h49;
s_mem_contents[14'h199c] = 8'hc3;
s_mem_contents[14'h199d] = 8'hc5;
s_mem_contents[14'h199e] = 8'h0c;
s_mem_contents[14'h199f] = 8'hd0;
s_mem_contents[14'h19a0] = 8'hfe;
s_mem_contents[14'h19a1] = 8'h68;
s_mem_contents[14'h19a2] = 8'h49;
s_mem_contents[14'h19a3] = 8'h30;
s_mem_contents[14'h19a4] = 8'hcd;
s_mem_contents[14'h19a5] = 8'h1f;
s_mem_contents[14'h19a6] = 8'h02;
s_mem_contents[14'h19a7] = 8'hd0;
s_mem_contents[14'h19a8] = 8'hfe;
s_mem_contents[14'h19a9] = 8'ha9;
s_mem_contents[14'h19aa] = 8'hff;
s_mem_contents[14'h19ab] = 8'h48;
s_mem_contents[14'h19ac] = 8'h28;
s_mem_contents[14'h19ad] = 8'had;
s_mem_contents[14'h19ae] = 8'h17;
s_mem_contents[14'h19af] = 8'h02;
s_mem_contents[14'h19b0] = 8'h08;
s_mem_contents[14'h19b1] = 8'h49;
s_mem_contents[14'h19b2] = 8'hc3;
s_mem_contents[14'h19b3] = 8'h28;
s_mem_contents[14'h19b4] = 8'h85;
s_mem_contents[14'h19b5] = 8'h02;
s_mem_contents[14'h19b6] = 8'h08;
s_mem_contents[14'h19b7] = 8'h49;
s_mem_contents[14'h19b8] = 8'hc3;
s_mem_contents[14'h19b9] = 8'hc5;
s_mem_contents[14'h19ba] = 8'h09;
s_mem_contents[14'h19bb] = 8'hd0;
s_mem_contents[14'h19bc] = 8'hfe;
s_mem_contents[14'h19bd] = 8'h68;
s_mem_contents[14'h19be] = 8'h49;
s_mem_contents[14'h19bf] = 8'h7d;
s_mem_contents[14'h19c0] = 8'hcd;
s_mem_contents[14'h19c1] = 8'h1c;
s_mem_contents[14'h19c2] = 8'h02;
s_mem_contents[14'h19c3] = 8'hd0;
s_mem_contents[14'h19c4] = 8'hfe;
s_mem_contents[14'h19c5] = 8'ha9;
s_mem_contents[14'h19c6] = 8'hff;
s_mem_contents[14'h19c7] = 8'h48;
s_mem_contents[14'h19c8] = 8'h28;
s_mem_contents[14'h19c9] = 8'had;
s_mem_contents[14'h19ca] = 8'h18;
s_mem_contents[14'h19cb] = 8'h02;
s_mem_contents[14'h19cc] = 8'h08;
s_mem_contents[14'h19cd] = 8'h49;
s_mem_contents[14'h19ce] = 8'hc3;
s_mem_contents[14'h19cf] = 8'h28;
s_mem_contents[14'h19d0] = 8'h85;
s_mem_contents[14'h19d1] = 8'h03;
s_mem_contents[14'h19d2] = 8'h08;
s_mem_contents[14'h19d3] = 8'h49;
s_mem_contents[14'h19d4] = 8'hc3;
s_mem_contents[14'h19d5] = 8'hc5;
s_mem_contents[14'h19d6] = 8'h0a;
s_mem_contents[14'h19d7] = 8'hd0;
s_mem_contents[14'h19d8] = 8'hfe;
s_mem_contents[14'h19d9] = 8'h68;
s_mem_contents[14'h19da] = 8'h49;
s_mem_contents[14'h19db] = 8'h7d;
s_mem_contents[14'h19dc] = 8'hcd;
s_mem_contents[14'h19dd] = 8'h1d;
s_mem_contents[14'h19de] = 8'h02;
s_mem_contents[14'h19df] = 8'hd0;
s_mem_contents[14'h19e0] = 8'hfe;
s_mem_contents[14'h19e1] = 8'ha9;
s_mem_contents[14'h19e2] = 8'hff;
s_mem_contents[14'h19e3] = 8'h48;
s_mem_contents[14'h19e4] = 8'h28;
s_mem_contents[14'h19e5] = 8'had;
s_mem_contents[14'h19e6] = 8'h19;
s_mem_contents[14'h19e7] = 8'h02;
s_mem_contents[14'h19e8] = 8'h08;
s_mem_contents[14'h19e9] = 8'h49;
s_mem_contents[14'h19ea] = 8'hc3;
s_mem_contents[14'h19eb] = 8'h28;
s_mem_contents[14'h19ec] = 8'h85;
s_mem_contents[14'h19ed] = 8'h04;
s_mem_contents[14'h19ee] = 8'h08;
s_mem_contents[14'h19ef] = 8'h49;
s_mem_contents[14'h19f0] = 8'hc3;
s_mem_contents[14'h19f1] = 8'hc5;
s_mem_contents[14'h19f2] = 8'h0b;
s_mem_contents[14'h19f3] = 8'hd0;
s_mem_contents[14'h19f4] = 8'hfe;
s_mem_contents[14'h19f5] = 8'h68;
s_mem_contents[14'h19f6] = 8'h49;
s_mem_contents[14'h19f7] = 8'h7d;
s_mem_contents[14'h19f8] = 8'hcd;
s_mem_contents[14'h19f9] = 8'h1e;
s_mem_contents[14'h19fa] = 8'h02;
s_mem_contents[14'h19fb] = 8'hd0;
s_mem_contents[14'h19fc] = 8'hfe;
s_mem_contents[14'h19fd] = 8'ha9;
s_mem_contents[14'h19fe] = 8'hff;
s_mem_contents[14'h19ff] = 8'h48;
s_mem_contents[14'h1a00] = 8'h28;
s_mem_contents[14'h1a01] = 8'had;
s_mem_contents[14'h1a02] = 8'h1a;
s_mem_contents[14'h1a03] = 8'h02;
s_mem_contents[14'h1a04] = 8'h08;
s_mem_contents[14'h1a05] = 8'h49;
s_mem_contents[14'h1a06] = 8'hc3;
s_mem_contents[14'h1a07] = 8'h28;
s_mem_contents[14'h1a08] = 8'h85;
s_mem_contents[14'h1a09] = 8'h05;
s_mem_contents[14'h1a0a] = 8'h08;
s_mem_contents[14'h1a0b] = 8'h49;
s_mem_contents[14'h1a0c] = 8'hc3;
s_mem_contents[14'h1a0d] = 8'hc5;
s_mem_contents[14'h1a0e] = 8'h0c;
s_mem_contents[14'h1a0f] = 8'hd0;
s_mem_contents[14'h1a10] = 8'hfe;
s_mem_contents[14'h1a11] = 8'h68;
s_mem_contents[14'h1a12] = 8'h49;
s_mem_contents[14'h1a13] = 8'h7d;
s_mem_contents[14'h1a14] = 8'hcd;
s_mem_contents[14'h1a15] = 8'h1f;
s_mem_contents[14'h1a16] = 8'h02;
s_mem_contents[14'h1a17] = 8'hd0;
s_mem_contents[14'h1a18] = 8'hfe;
s_mem_contents[14'h1a19] = 8'ha9;
s_mem_contents[14'h1a1a] = 8'h00;
s_mem_contents[14'h1a1b] = 8'h48;
s_mem_contents[14'h1a1c] = 8'h28;
s_mem_contents[14'h1a1d] = 8'ha9;
s_mem_contents[14'h1a1e] = 8'hc3;
s_mem_contents[14'h1a1f] = 8'h08;
s_mem_contents[14'h1a20] = 8'hcd;
s_mem_contents[14'h1a21] = 8'h17;
s_mem_contents[14'h1a22] = 8'h02;
s_mem_contents[14'h1a23] = 8'hd0;
s_mem_contents[14'h1a24] = 8'hfe;
s_mem_contents[14'h1a25] = 8'h68;
s_mem_contents[14'h1a26] = 8'h49;
s_mem_contents[14'h1a27] = 8'h30;
s_mem_contents[14'h1a28] = 8'hcd;
s_mem_contents[14'h1a29] = 8'h1c;
s_mem_contents[14'h1a2a] = 8'h02;
s_mem_contents[14'h1a2b] = 8'hd0;
s_mem_contents[14'h1a2c] = 8'hfe;
s_mem_contents[14'h1a2d] = 8'ha9;
s_mem_contents[14'h1a2e] = 8'h00;
s_mem_contents[14'h1a2f] = 8'h48;
s_mem_contents[14'h1a30] = 8'h28;
s_mem_contents[14'h1a31] = 8'ha9;
s_mem_contents[14'h1a32] = 8'h82;
s_mem_contents[14'h1a33] = 8'h08;
s_mem_contents[14'h1a34] = 8'hcd;
s_mem_contents[14'h1a35] = 8'h18;
s_mem_contents[14'h1a36] = 8'h02;
s_mem_contents[14'h1a37] = 8'hd0;
s_mem_contents[14'h1a38] = 8'hfe;
s_mem_contents[14'h1a39] = 8'h68;
s_mem_contents[14'h1a3a] = 8'h49;
s_mem_contents[14'h1a3b] = 8'h30;
s_mem_contents[14'h1a3c] = 8'hcd;
s_mem_contents[14'h1a3d] = 8'h1d;
s_mem_contents[14'h1a3e] = 8'h02;
s_mem_contents[14'h1a3f] = 8'hd0;
s_mem_contents[14'h1a40] = 8'hfe;
s_mem_contents[14'h1a41] = 8'ha9;
s_mem_contents[14'h1a42] = 8'h00;
s_mem_contents[14'h1a43] = 8'h48;
s_mem_contents[14'h1a44] = 8'h28;
s_mem_contents[14'h1a45] = 8'ha9;
s_mem_contents[14'h1a46] = 8'h41;
s_mem_contents[14'h1a47] = 8'h08;
s_mem_contents[14'h1a48] = 8'hcd;
s_mem_contents[14'h1a49] = 8'h19;
s_mem_contents[14'h1a4a] = 8'h02;
s_mem_contents[14'h1a4b] = 8'hd0;
s_mem_contents[14'h1a4c] = 8'hfe;
s_mem_contents[14'h1a4d] = 8'h68;
s_mem_contents[14'h1a4e] = 8'h49;
s_mem_contents[14'h1a4f] = 8'h30;
s_mem_contents[14'h1a50] = 8'hcd;
s_mem_contents[14'h1a51] = 8'h1e;
s_mem_contents[14'h1a52] = 8'h02;
s_mem_contents[14'h1a53] = 8'hd0;
s_mem_contents[14'h1a54] = 8'hfe;
s_mem_contents[14'h1a55] = 8'ha9;
s_mem_contents[14'h1a56] = 8'h00;
s_mem_contents[14'h1a57] = 8'h48;
s_mem_contents[14'h1a58] = 8'h28;
s_mem_contents[14'h1a59] = 8'ha9;
s_mem_contents[14'h1a5a] = 8'h00;
s_mem_contents[14'h1a5b] = 8'h08;
s_mem_contents[14'h1a5c] = 8'hcd;
s_mem_contents[14'h1a5d] = 8'h1a;
s_mem_contents[14'h1a5e] = 8'h02;
s_mem_contents[14'h1a5f] = 8'hd0;
s_mem_contents[14'h1a60] = 8'hfe;
s_mem_contents[14'h1a61] = 8'h68;
s_mem_contents[14'h1a62] = 8'h49;
s_mem_contents[14'h1a63] = 8'h30;
s_mem_contents[14'h1a64] = 8'hcd;
s_mem_contents[14'h1a65] = 8'h1f;
s_mem_contents[14'h1a66] = 8'h02;
s_mem_contents[14'h1a67] = 8'hd0;
s_mem_contents[14'h1a68] = 8'hfe;
s_mem_contents[14'h1a69] = 8'ha9;
s_mem_contents[14'h1a6a] = 8'hff;
s_mem_contents[14'h1a6b] = 8'h48;
s_mem_contents[14'h1a6c] = 8'h28;
s_mem_contents[14'h1a6d] = 8'ha9;
s_mem_contents[14'h1a6e] = 8'hc3;
s_mem_contents[14'h1a6f] = 8'h08;
s_mem_contents[14'h1a70] = 8'hcd;
s_mem_contents[14'h1a71] = 8'h17;
s_mem_contents[14'h1a72] = 8'h02;
s_mem_contents[14'h1a73] = 8'hd0;
s_mem_contents[14'h1a74] = 8'hfe;
s_mem_contents[14'h1a75] = 8'h68;
s_mem_contents[14'h1a76] = 8'h49;
s_mem_contents[14'h1a77] = 8'h7d;
s_mem_contents[14'h1a78] = 8'hcd;
s_mem_contents[14'h1a79] = 8'h1c;
s_mem_contents[14'h1a7a] = 8'h02;
s_mem_contents[14'h1a7b] = 8'hd0;
s_mem_contents[14'h1a7c] = 8'hfe;
s_mem_contents[14'h1a7d] = 8'ha9;
s_mem_contents[14'h1a7e] = 8'hff;
s_mem_contents[14'h1a7f] = 8'h48;
s_mem_contents[14'h1a80] = 8'h28;
s_mem_contents[14'h1a81] = 8'ha9;
s_mem_contents[14'h1a82] = 8'h82;
s_mem_contents[14'h1a83] = 8'h08;
s_mem_contents[14'h1a84] = 8'hcd;
s_mem_contents[14'h1a85] = 8'h18;
s_mem_contents[14'h1a86] = 8'h02;
s_mem_contents[14'h1a87] = 8'hd0;
s_mem_contents[14'h1a88] = 8'hfe;
s_mem_contents[14'h1a89] = 8'h68;
s_mem_contents[14'h1a8a] = 8'h49;
s_mem_contents[14'h1a8b] = 8'h7d;
s_mem_contents[14'h1a8c] = 8'hcd;
s_mem_contents[14'h1a8d] = 8'h1d;
s_mem_contents[14'h1a8e] = 8'h02;
s_mem_contents[14'h1a8f] = 8'hd0;
s_mem_contents[14'h1a90] = 8'hfe;
s_mem_contents[14'h1a91] = 8'ha9;
s_mem_contents[14'h1a92] = 8'hff;
s_mem_contents[14'h1a93] = 8'h48;
s_mem_contents[14'h1a94] = 8'h28;
s_mem_contents[14'h1a95] = 8'ha9;
s_mem_contents[14'h1a96] = 8'h41;
s_mem_contents[14'h1a97] = 8'h08;
s_mem_contents[14'h1a98] = 8'hcd;
s_mem_contents[14'h1a99] = 8'h19;
s_mem_contents[14'h1a9a] = 8'h02;
s_mem_contents[14'h1a9b] = 8'hd0;
s_mem_contents[14'h1a9c] = 8'hfe;
s_mem_contents[14'h1a9d] = 8'h68;
s_mem_contents[14'h1a9e] = 8'h49;
s_mem_contents[14'h1a9f] = 8'h7d;
s_mem_contents[14'h1aa0] = 8'hcd;
s_mem_contents[14'h1aa1] = 8'h1e;
s_mem_contents[14'h1aa2] = 8'h02;
s_mem_contents[14'h1aa3] = 8'hd0;
s_mem_contents[14'h1aa4] = 8'hfe;
s_mem_contents[14'h1aa5] = 8'ha9;
s_mem_contents[14'h1aa6] = 8'hff;
s_mem_contents[14'h1aa7] = 8'h48;
s_mem_contents[14'h1aa8] = 8'h28;
s_mem_contents[14'h1aa9] = 8'ha9;
s_mem_contents[14'h1aaa] = 8'h00;
s_mem_contents[14'h1aab] = 8'h08;
s_mem_contents[14'h1aac] = 8'hcd;
s_mem_contents[14'h1aad] = 8'h1a;
s_mem_contents[14'h1aae] = 8'h02;
s_mem_contents[14'h1aaf] = 8'hd0;
s_mem_contents[14'h1ab0] = 8'hfe;
s_mem_contents[14'h1ab1] = 8'h68;
s_mem_contents[14'h1ab2] = 8'h49;
s_mem_contents[14'h1ab3] = 8'h7d;
s_mem_contents[14'h1ab4] = 8'hcd;
s_mem_contents[14'h1ab5] = 8'h1f;
s_mem_contents[14'h1ab6] = 8'h02;
s_mem_contents[14'h1ab7] = 8'hd0;
s_mem_contents[14'h1ab8] = 8'hfe;
s_mem_contents[14'h1ab9] = 8'ha2;
s_mem_contents[14'h1aba] = 8'h00;
s_mem_contents[14'h1abb] = 8'ha5;
s_mem_contents[14'h1abc] = 8'h02;
s_mem_contents[14'h1abd] = 8'h49;
s_mem_contents[14'h1abe] = 8'hc3;
s_mem_contents[14'h1abf] = 8'hc5;
s_mem_contents[14'h1ac0] = 8'h09;
s_mem_contents[14'h1ac1] = 8'hd0;
s_mem_contents[14'h1ac2] = 8'hfe;
s_mem_contents[14'h1ac3] = 8'h86;
s_mem_contents[14'h1ac4] = 8'h02;
s_mem_contents[14'h1ac5] = 8'had;
s_mem_contents[14'h1ac6] = 8'h03;
s_mem_contents[14'h1ac7] = 8'h02;
s_mem_contents[14'h1ac8] = 8'h49;
s_mem_contents[14'h1ac9] = 8'hc3;
s_mem_contents[14'h1aca] = 8'hcd;
s_mem_contents[14'h1acb] = 8'h17;
s_mem_contents[14'h1acc] = 8'h02;
s_mem_contents[14'h1acd] = 8'hd0;
s_mem_contents[14'h1ace] = 8'hfe;
s_mem_contents[14'h1acf] = 8'h8e;
s_mem_contents[14'h1ad0] = 8'h03;
s_mem_contents[14'h1ad1] = 8'h02;
s_mem_contents[14'h1ad2] = 8'ha5;
s_mem_contents[14'h1ad3] = 8'h03;
s_mem_contents[14'h1ad4] = 8'h49;
s_mem_contents[14'h1ad5] = 8'hc3;
s_mem_contents[14'h1ad6] = 8'hc5;
s_mem_contents[14'h1ad7] = 8'h0a;
s_mem_contents[14'h1ad8] = 8'hd0;
s_mem_contents[14'h1ad9] = 8'hfe;
s_mem_contents[14'h1ada] = 8'h86;
s_mem_contents[14'h1adb] = 8'h03;
s_mem_contents[14'h1adc] = 8'had;
s_mem_contents[14'h1add] = 8'h04;
s_mem_contents[14'h1ade] = 8'h02;
s_mem_contents[14'h1adf] = 8'h49;
s_mem_contents[14'h1ae0] = 8'hc3;
s_mem_contents[14'h1ae1] = 8'hcd;
s_mem_contents[14'h1ae2] = 8'h18;
s_mem_contents[14'h1ae3] = 8'h02;
s_mem_contents[14'h1ae4] = 8'hd0;
s_mem_contents[14'h1ae5] = 8'hfe;
s_mem_contents[14'h1ae6] = 8'h8e;
s_mem_contents[14'h1ae7] = 8'h04;
s_mem_contents[14'h1ae8] = 8'h02;
s_mem_contents[14'h1ae9] = 8'ha5;
s_mem_contents[14'h1aea] = 8'h04;
s_mem_contents[14'h1aeb] = 8'h49;
s_mem_contents[14'h1aec] = 8'hc3;
s_mem_contents[14'h1aed] = 8'hc5;
s_mem_contents[14'h1aee] = 8'h0b;
s_mem_contents[14'h1aef] = 8'hd0;
s_mem_contents[14'h1af0] = 8'hfe;
s_mem_contents[14'h1af1] = 8'h86;
s_mem_contents[14'h1af2] = 8'h04;
s_mem_contents[14'h1af3] = 8'had;
s_mem_contents[14'h1af4] = 8'h05;
s_mem_contents[14'h1af5] = 8'h02;
s_mem_contents[14'h1af6] = 8'h49;
s_mem_contents[14'h1af7] = 8'hc3;
s_mem_contents[14'h1af8] = 8'hcd;
s_mem_contents[14'h1af9] = 8'h19;
s_mem_contents[14'h1afa] = 8'h02;
s_mem_contents[14'h1afb] = 8'hd0;
s_mem_contents[14'h1afc] = 8'hfe;
s_mem_contents[14'h1afd] = 8'h8e;
s_mem_contents[14'h1afe] = 8'h05;
s_mem_contents[14'h1aff] = 8'h02;
s_mem_contents[14'h1b00] = 8'ha5;
s_mem_contents[14'h1b01] = 8'h05;
s_mem_contents[14'h1b02] = 8'h49;
s_mem_contents[14'h1b03] = 8'hc3;
s_mem_contents[14'h1b04] = 8'hc5;
s_mem_contents[14'h1b05] = 8'h0c;
s_mem_contents[14'h1b06] = 8'hd0;
s_mem_contents[14'h1b07] = 8'hfe;
s_mem_contents[14'h1b08] = 8'h86;
s_mem_contents[14'h1b09] = 8'h05;
s_mem_contents[14'h1b0a] = 8'had;
s_mem_contents[14'h1b0b] = 8'h06;
s_mem_contents[14'h1b0c] = 8'h02;
s_mem_contents[14'h1b0d] = 8'h49;
s_mem_contents[14'h1b0e] = 8'hc3;
s_mem_contents[14'h1b0f] = 8'hcd;
s_mem_contents[14'h1b10] = 8'h1a;
s_mem_contents[14'h1b11] = 8'h02;
s_mem_contents[14'h1b12] = 8'hd0;
s_mem_contents[14'h1b13] = 8'hfe;
s_mem_contents[14'h1b14] = 8'h8e;
s_mem_contents[14'h1b15] = 8'h06;
s_mem_contents[14'h1b16] = 8'h02;
s_mem_contents[14'h1b17] = 8'had;
s_mem_contents[14'h1b18] = 8'h00;
s_mem_contents[14'h1b19] = 8'h02;
s_mem_contents[14'h1b1a] = 8'hc9;
s_mem_contents[14'h1b1b] = 8'h18;
s_mem_contents[14'h1b1c] = 8'hd0;
s_mem_contents[14'h1b1d] = 8'hfe;
s_mem_contents[14'h1b1e] = 8'ha9;
s_mem_contents[14'h1b1f] = 8'h19;
s_mem_contents[14'h1b20] = 8'h8d;
s_mem_contents[14'h1b21] = 8'h00;
s_mem_contents[14'h1b22] = 8'h02;
s_mem_contents[14'h1b23] = 8'ha9;
s_mem_contents[14'h1b24] = 8'h00;
s_mem_contents[14'h1b25] = 8'h48;
s_mem_contents[14'h1b26] = 8'ha9;
s_mem_contents[14'h1b27] = 8'hff;
s_mem_contents[14'h1b28] = 8'h28;
s_mem_contents[14'h1b29] = 8'h24;
s_mem_contents[14'h1b2a] = 8'h0c;
s_mem_contents[14'h1b2b] = 8'h08;
s_mem_contents[14'h1b2c] = 8'hc9;
s_mem_contents[14'h1b2d] = 8'hff;
s_mem_contents[14'h1b2e] = 8'hd0;
s_mem_contents[14'h1b2f] = 8'hfe;
s_mem_contents[14'h1b30] = 8'h68;
s_mem_contents[14'h1b31] = 8'h48;
s_mem_contents[14'h1b32] = 8'hc9;
s_mem_contents[14'h1b33] = 8'h32;
s_mem_contents[14'h1b34] = 8'hd0;
s_mem_contents[14'h1b35] = 8'hfe;
s_mem_contents[14'h1b36] = 8'h28;
s_mem_contents[14'h1b37] = 8'ha9;
s_mem_contents[14'h1b38] = 8'h00;
s_mem_contents[14'h1b39] = 8'h48;
s_mem_contents[14'h1b3a] = 8'ha9;
s_mem_contents[14'h1b3b] = 8'h01;
s_mem_contents[14'h1b3c] = 8'h28;
s_mem_contents[14'h1b3d] = 8'h24;
s_mem_contents[14'h1b3e] = 8'h0b;
s_mem_contents[14'h1b3f] = 8'h08;
s_mem_contents[14'h1b40] = 8'hc9;
s_mem_contents[14'h1b41] = 8'h01;
s_mem_contents[14'h1b42] = 8'hd0;
s_mem_contents[14'h1b43] = 8'hfe;
s_mem_contents[14'h1b44] = 8'h68;
s_mem_contents[14'h1b45] = 8'h48;
s_mem_contents[14'h1b46] = 8'hc9;
s_mem_contents[14'h1b47] = 8'h70;
s_mem_contents[14'h1b48] = 8'hd0;
s_mem_contents[14'h1b49] = 8'hfe;
s_mem_contents[14'h1b4a] = 8'h28;
s_mem_contents[14'h1b4b] = 8'ha9;
s_mem_contents[14'h1b4c] = 8'h00;
s_mem_contents[14'h1b4d] = 8'h48;
s_mem_contents[14'h1b4e] = 8'ha9;
s_mem_contents[14'h1b4f] = 8'h01;
s_mem_contents[14'h1b50] = 8'h28;
s_mem_contents[14'h1b51] = 8'h24;
s_mem_contents[14'h1b52] = 8'h0a;
s_mem_contents[14'h1b53] = 8'h08;
s_mem_contents[14'h1b54] = 8'hc9;
s_mem_contents[14'h1b55] = 8'h01;
s_mem_contents[14'h1b56] = 8'hd0;
s_mem_contents[14'h1b57] = 8'hfe;
s_mem_contents[14'h1b58] = 8'h68;
s_mem_contents[14'h1b59] = 8'h48;
s_mem_contents[14'h1b5a] = 8'hc9;
s_mem_contents[14'h1b5b] = 8'hb2;
s_mem_contents[14'h1b5c] = 8'hd0;
s_mem_contents[14'h1b5d] = 8'hfe;
s_mem_contents[14'h1b5e] = 8'h28;
s_mem_contents[14'h1b5f] = 8'ha9;
s_mem_contents[14'h1b60] = 8'h00;
s_mem_contents[14'h1b61] = 8'h48;
s_mem_contents[14'h1b62] = 8'ha9;
s_mem_contents[14'h1b63] = 8'h01;
s_mem_contents[14'h1b64] = 8'h28;
s_mem_contents[14'h1b65] = 8'h24;
s_mem_contents[14'h1b66] = 8'h09;
s_mem_contents[14'h1b67] = 8'h08;
s_mem_contents[14'h1b68] = 8'hc9;
s_mem_contents[14'h1b69] = 8'h01;
s_mem_contents[14'h1b6a] = 8'hd0;
s_mem_contents[14'h1b6b] = 8'hfe;
s_mem_contents[14'h1b6c] = 8'h68;
s_mem_contents[14'h1b6d] = 8'h48;
s_mem_contents[14'h1b6e] = 8'hc9;
s_mem_contents[14'h1b6f] = 8'hf0;
s_mem_contents[14'h1b70] = 8'hd0;
s_mem_contents[14'h1b71] = 8'hfe;
s_mem_contents[14'h1b72] = 8'h28;
s_mem_contents[14'h1b73] = 8'ha9;
s_mem_contents[14'h1b74] = 8'hff;
s_mem_contents[14'h1b75] = 8'h48;
s_mem_contents[14'h1b76] = 8'ha9;
s_mem_contents[14'h1b77] = 8'hff;
s_mem_contents[14'h1b78] = 8'h28;
s_mem_contents[14'h1b79] = 8'h24;
s_mem_contents[14'h1b7a] = 8'h0c;
s_mem_contents[14'h1b7b] = 8'h08;
s_mem_contents[14'h1b7c] = 8'hc9;
s_mem_contents[14'h1b7d] = 8'hff;
s_mem_contents[14'h1b7e] = 8'hd0;
s_mem_contents[14'h1b7f] = 8'hfe;
s_mem_contents[14'h1b80] = 8'h68;
s_mem_contents[14'h1b81] = 8'h48;
s_mem_contents[14'h1b82] = 8'hc9;
s_mem_contents[14'h1b83] = 8'h3f;
s_mem_contents[14'h1b84] = 8'hd0;
s_mem_contents[14'h1b85] = 8'hfe;
s_mem_contents[14'h1b86] = 8'h28;
s_mem_contents[14'h1b87] = 8'ha9;
s_mem_contents[14'h1b88] = 8'hff;
s_mem_contents[14'h1b89] = 8'h48;
s_mem_contents[14'h1b8a] = 8'ha9;
s_mem_contents[14'h1b8b] = 8'h01;
s_mem_contents[14'h1b8c] = 8'h28;
s_mem_contents[14'h1b8d] = 8'h24;
s_mem_contents[14'h1b8e] = 8'h0b;
s_mem_contents[14'h1b8f] = 8'h08;
s_mem_contents[14'h1b90] = 8'hc9;
s_mem_contents[14'h1b91] = 8'h01;
s_mem_contents[14'h1b92] = 8'hd0;
s_mem_contents[14'h1b93] = 8'hfe;
s_mem_contents[14'h1b94] = 8'h68;
s_mem_contents[14'h1b95] = 8'h48;
s_mem_contents[14'h1b96] = 8'hc9;
s_mem_contents[14'h1b97] = 8'h7d;
s_mem_contents[14'h1b98] = 8'hd0;
s_mem_contents[14'h1b99] = 8'hfe;
s_mem_contents[14'h1b9a] = 8'h28;
s_mem_contents[14'h1b9b] = 8'ha9;
s_mem_contents[14'h1b9c] = 8'hff;
s_mem_contents[14'h1b9d] = 8'h48;
s_mem_contents[14'h1b9e] = 8'ha9;
s_mem_contents[14'h1b9f] = 8'h01;
s_mem_contents[14'h1ba0] = 8'h28;
s_mem_contents[14'h1ba1] = 8'h24;
s_mem_contents[14'h1ba2] = 8'h0a;
s_mem_contents[14'h1ba3] = 8'h08;
s_mem_contents[14'h1ba4] = 8'hc9;
s_mem_contents[14'h1ba5] = 8'h01;
s_mem_contents[14'h1ba6] = 8'hd0;
s_mem_contents[14'h1ba7] = 8'hfe;
s_mem_contents[14'h1ba8] = 8'h68;
s_mem_contents[14'h1ba9] = 8'h48;
s_mem_contents[14'h1baa] = 8'hc9;
s_mem_contents[14'h1bab] = 8'hbf;
s_mem_contents[14'h1bac] = 8'hd0;
s_mem_contents[14'h1bad] = 8'hfe;
s_mem_contents[14'h1bae] = 8'h28;
s_mem_contents[14'h1baf] = 8'ha9;
s_mem_contents[14'h1bb0] = 8'hff;
s_mem_contents[14'h1bb1] = 8'h48;
s_mem_contents[14'h1bb2] = 8'ha9;
s_mem_contents[14'h1bb3] = 8'h01;
s_mem_contents[14'h1bb4] = 8'h28;
s_mem_contents[14'h1bb5] = 8'h24;
s_mem_contents[14'h1bb6] = 8'h09;
s_mem_contents[14'h1bb7] = 8'h08;
s_mem_contents[14'h1bb8] = 8'hc9;
s_mem_contents[14'h1bb9] = 8'h01;
s_mem_contents[14'h1bba] = 8'hd0;
s_mem_contents[14'h1bbb] = 8'hfe;
s_mem_contents[14'h1bbc] = 8'h68;
s_mem_contents[14'h1bbd] = 8'h48;
s_mem_contents[14'h1bbe] = 8'hc9;
s_mem_contents[14'h1bbf] = 8'hfd;
s_mem_contents[14'h1bc0] = 8'hd0;
s_mem_contents[14'h1bc1] = 8'hfe;
s_mem_contents[14'h1bc2] = 8'h28;
s_mem_contents[14'h1bc3] = 8'ha9;
s_mem_contents[14'h1bc4] = 8'h00;
s_mem_contents[14'h1bc5] = 8'h48;
s_mem_contents[14'h1bc6] = 8'ha9;
s_mem_contents[14'h1bc7] = 8'hff;
s_mem_contents[14'h1bc8] = 8'h28;
s_mem_contents[14'h1bc9] = 8'h2c;
s_mem_contents[14'h1bca] = 8'h1a;
s_mem_contents[14'h1bcb] = 8'h02;
s_mem_contents[14'h1bcc] = 8'h08;
s_mem_contents[14'h1bcd] = 8'hc9;
s_mem_contents[14'h1bce] = 8'hff;
s_mem_contents[14'h1bcf] = 8'hd0;
s_mem_contents[14'h1bd0] = 8'hfe;
s_mem_contents[14'h1bd1] = 8'h68;
s_mem_contents[14'h1bd2] = 8'h48;
s_mem_contents[14'h1bd3] = 8'hc9;
s_mem_contents[14'h1bd4] = 8'h32;
s_mem_contents[14'h1bd5] = 8'hd0;
s_mem_contents[14'h1bd6] = 8'hfe;
s_mem_contents[14'h1bd7] = 8'h28;
s_mem_contents[14'h1bd8] = 8'ha9;
s_mem_contents[14'h1bd9] = 8'h00;
s_mem_contents[14'h1bda] = 8'h48;
s_mem_contents[14'h1bdb] = 8'ha9;
s_mem_contents[14'h1bdc] = 8'h01;
s_mem_contents[14'h1bdd] = 8'h28;
s_mem_contents[14'h1bde] = 8'h2c;
s_mem_contents[14'h1bdf] = 8'h19;
s_mem_contents[14'h1be0] = 8'h02;
s_mem_contents[14'h1be1] = 8'h08;
s_mem_contents[14'h1be2] = 8'hc9;
s_mem_contents[14'h1be3] = 8'h01;
s_mem_contents[14'h1be4] = 8'hd0;
s_mem_contents[14'h1be5] = 8'hfe;
s_mem_contents[14'h1be6] = 8'h68;
s_mem_contents[14'h1be7] = 8'h48;
s_mem_contents[14'h1be8] = 8'hc9;
s_mem_contents[14'h1be9] = 8'h70;
s_mem_contents[14'h1bea] = 8'hd0;
s_mem_contents[14'h1beb] = 8'hfe;
s_mem_contents[14'h1bec] = 8'h28;
s_mem_contents[14'h1bed] = 8'ha9;
s_mem_contents[14'h1bee] = 8'h00;
s_mem_contents[14'h1bef] = 8'h48;
s_mem_contents[14'h1bf0] = 8'ha9;
s_mem_contents[14'h1bf1] = 8'h01;
s_mem_contents[14'h1bf2] = 8'h28;
s_mem_contents[14'h1bf3] = 8'h2c;
s_mem_contents[14'h1bf4] = 8'h18;
s_mem_contents[14'h1bf5] = 8'h02;
s_mem_contents[14'h1bf6] = 8'h08;
s_mem_contents[14'h1bf7] = 8'hc9;
s_mem_contents[14'h1bf8] = 8'h01;
s_mem_contents[14'h1bf9] = 8'hd0;
s_mem_contents[14'h1bfa] = 8'hfe;
s_mem_contents[14'h1bfb] = 8'h68;
s_mem_contents[14'h1bfc] = 8'h48;
s_mem_contents[14'h1bfd] = 8'hc9;
s_mem_contents[14'h1bfe] = 8'hb2;
s_mem_contents[14'h1bff] = 8'hd0;
s_mem_contents[14'h1c00] = 8'hfe;
s_mem_contents[14'h1c01] = 8'h28;
s_mem_contents[14'h1c02] = 8'ha9;
s_mem_contents[14'h1c03] = 8'h00;
s_mem_contents[14'h1c04] = 8'h48;
s_mem_contents[14'h1c05] = 8'ha9;
s_mem_contents[14'h1c06] = 8'h01;
s_mem_contents[14'h1c07] = 8'h28;
s_mem_contents[14'h1c08] = 8'h2c;
s_mem_contents[14'h1c09] = 8'h17;
s_mem_contents[14'h1c0a] = 8'h02;
s_mem_contents[14'h1c0b] = 8'h08;
s_mem_contents[14'h1c0c] = 8'hc9;
s_mem_contents[14'h1c0d] = 8'h01;
s_mem_contents[14'h1c0e] = 8'hd0;
s_mem_contents[14'h1c0f] = 8'hfe;
s_mem_contents[14'h1c10] = 8'h68;
s_mem_contents[14'h1c11] = 8'h48;
s_mem_contents[14'h1c12] = 8'hc9;
s_mem_contents[14'h1c13] = 8'hf0;
s_mem_contents[14'h1c14] = 8'hd0;
s_mem_contents[14'h1c15] = 8'hfe;
s_mem_contents[14'h1c16] = 8'h28;
s_mem_contents[14'h1c17] = 8'ha9;
s_mem_contents[14'h1c18] = 8'hff;
s_mem_contents[14'h1c19] = 8'h48;
s_mem_contents[14'h1c1a] = 8'ha9;
s_mem_contents[14'h1c1b] = 8'hff;
s_mem_contents[14'h1c1c] = 8'h28;
s_mem_contents[14'h1c1d] = 8'h2c;
s_mem_contents[14'h1c1e] = 8'h1a;
s_mem_contents[14'h1c1f] = 8'h02;
s_mem_contents[14'h1c20] = 8'h08;
s_mem_contents[14'h1c21] = 8'hc9;
s_mem_contents[14'h1c22] = 8'hff;
s_mem_contents[14'h1c23] = 8'hd0;
s_mem_contents[14'h1c24] = 8'hfe;
s_mem_contents[14'h1c25] = 8'h68;
s_mem_contents[14'h1c26] = 8'h48;
s_mem_contents[14'h1c27] = 8'hc9;
s_mem_contents[14'h1c28] = 8'h3f;
s_mem_contents[14'h1c29] = 8'hd0;
s_mem_contents[14'h1c2a] = 8'hfe;
s_mem_contents[14'h1c2b] = 8'h28;
s_mem_contents[14'h1c2c] = 8'ha9;
s_mem_contents[14'h1c2d] = 8'hff;
s_mem_contents[14'h1c2e] = 8'h48;
s_mem_contents[14'h1c2f] = 8'ha9;
s_mem_contents[14'h1c30] = 8'h01;
s_mem_contents[14'h1c31] = 8'h28;
s_mem_contents[14'h1c32] = 8'h2c;
s_mem_contents[14'h1c33] = 8'h19;
s_mem_contents[14'h1c34] = 8'h02;
s_mem_contents[14'h1c35] = 8'h08;
s_mem_contents[14'h1c36] = 8'hc9;
s_mem_contents[14'h1c37] = 8'h01;
s_mem_contents[14'h1c38] = 8'hd0;
s_mem_contents[14'h1c39] = 8'hfe;
s_mem_contents[14'h1c3a] = 8'h68;
s_mem_contents[14'h1c3b] = 8'h48;
s_mem_contents[14'h1c3c] = 8'hc9;
s_mem_contents[14'h1c3d] = 8'h7d;
s_mem_contents[14'h1c3e] = 8'hd0;
s_mem_contents[14'h1c3f] = 8'hfe;
s_mem_contents[14'h1c40] = 8'h28;
s_mem_contents[14'h1c41] = 8'ha9;
s_mem_contents[14'h1c42] = 8'hff;
s_mem_contents[14'h1c43] = 8'h48;
s_mem_contents[14'h1c44] = 8'ha9;
s_mem_contents[14'h1c45] = 8'h01;
s_mem_contents[14'h1c46] = 8'h28;
s_mem_contents[14'h1c47] = 8'h2c;
s_mem_contents[14'h1c48] = 8'h18;
s_mem_contents[14'h1c49] = 8'h02;
s_mem_contents[14'h1c4a] = 8'h08;
s_mem_contents[14'h1c4b] = 8'hc9;
s_mem_contents[14'h1c4c] = 8'h01;
s_mem_contents[14'h1c4d] = 8'hd0;
s_mem_contents[14'h1c4e] = 8'hfe;
s_mem_contents[14'h1c4f] = 8'h68;
s_mem_contents[14'h1c50] = 8'h48;
s_mem_contents[14'h1c51] = 8'hc9;
s_mem_contents[14'h1c52] = 8'hbf;
s_mem_contents[14'h1c53] = 8'hd0;
s_mem_contents[14'h1c54] = 8'hfe;
s_mem_contents[14'h1c55] = 8'h28;
s_mem_contents[14'h1c56] = 8'ha9;
s_mem_contents[14'h1c57] = 8'hff;
s_mem_contents[14'h1c58] = 8'h48;
s_mem_contents[14'h1c59] = 8'ha9;
s_mem_contents[14'h1c5a] = 8'h01;
s_mem_contents[14'h1c5b] = 8'h28;
s_mem_contents[14'h1c5c] = 8'h2c;
s_mem_contents[14'h1c5d] = 8'h17;
s_mem_contents[14'h1c5e] = 8'h02;
s_mem_contents[14'h1c5f] = 8'h08;
s_mem_contents[14'h1c60] = 8'hc9;
s_mem_contents[14'h1c61] = 8'h01;
s_mem_contents[14'h1c62] = 8'hd0;
s_mem_contents[14'h1c63] = 8'hfe;
s_mem_contents[14'h1c64] = 8'h68;
s_mem_contents[14'h1c65] = 8'h48;
s_mem_contents[14'h1c66] = 8'hc9;
s_mem_contents[14'h1c67] = 8'hfd;
s_mem_contents[14'h1c68] = 8'hd0;
s_mem_contents[14'h1c69] = 8'hfe;
s_mem_contents[14'h1c6a] = 8'h28;
s_mem_contents[14'h1c6b] = 8'had;
s_mem_contents[14'h1c6c] = 8'h00;
s_mem_contents[14'h1c6d] = 8'h02;
s_mem_contents[14'h1c6e] = 8'hc9;
s_mem_contents[14'h1c6f] = 8'h19;
s_mem_contents[14'h1c70] = 8'hd0;
s_mem_contents[14'h1c71] = 8'hfe;
s_mem_contents[14'h1c72] = 8'ha9;
s_mem_contents[14'h1c73] = 8'h1a;
s_mem_contents[14'h1c74] = 8'h8d;
s_mem_contents[14'h1c75] = 8'h00;
s_mem_contents[14'h1c76] = 8'h02;
s_mem_contents[14'h1c77] = 8'ha9;
s_mem_contents[14'h1c78] = 8'h00;
s_mem_contents[14'h1c79] = 8'h48;
s_mem_contents[14'h1c7a] = 8'ha2;
s_mem_contents[14'h1c7b] = 8'h80;
s_mem_contents[14'h1c7c] = 8'h28;
s_mem_contents[14'h1c7d] = 8'he4;
s_mem_contents[14'h1c7e] = 8'h0d;
s_mem_contents[14'h1c7f] = 8'h08;
s_mem_contents[14'h1c80] = 8'h68;
s_mem_contents[14'h1c81] = 8'h48;
s_mem_contents[14'h1c82] = 8'hc9;
s_mem_contents[14'h1c83] = 8'h31;
s_mem_contents[14'h1c84] = 8'hd0;
s_mem_contents[14'h1c85] = 8'hfe;
s_mem_contents[14'h1c86] = 8'h28;
s_mem_contents[14'h1c87] = 8'hca;
s_mem_contents[14'h1c88] = 8'he4;
s_mem_contents[14'h1c89] = 8'h0d;
s_mem_contents[14'h1c8a] = 8'h08;
s_mem_contents[14'h1c8b] = 8'h68;
s_mem_contents[14'h1c8c] = 8'h48;
s_mem_contents[14'h1c8d] = 8'hc9;
s_mem_contents[14'h1c8e] = 8'h33;
s_mem_contents[14'h1c8f] = 8'hd0;
s_mem_contents[14'h1c90] = 8'hfe;
s_mem_contents[14'h1c91] = 8'h28;
s_mem_contents[14'h1c92] = 8'hca;
s_mem_contents[14'h1c93] = 8'he4;
s_mem_contents[14'h1c94] = 8'h0d;
s_mem_contents[14'h1c95] = 8'h08;
s_mem_contents[14'h1c96] = 8'he0;
s_mem_contents[14'h1c97] = 8'h7e;
s_mem_contents[14'h1c98] = 8'hd0;
s_mem_contents[14'h1c99] = 8'hfe;
s_mem_contents[14'h1c9a] = 8'h68;
s_mem_contents[14'h1c9b] = 8'h48;
s_mem_contents[14'h1c9c] = 8'hc9;
s_mem_contents[14'h1c9d] = 8'hb0;
s_mem_contents[14'h1c9e] = 8'hd0;
s_mem_contents[14'h1c9f] = 8'hfe;
s_mem_contents[14'h1ca0] = 8'h28;
s_mem_contents[14'h1ca1] = 8'ha9;
s_mem_contents[14'h1ca2] = 8'hff;
s_mem_contents[14'h1ca3] = 8'h48;
s_mem_contents[14'h1ca4] = 8'ha2;
s_mem_contents[14'h1ca5] = 8'h80;
s_mem_contents[14'h1ca6] = 8'h28;
s_mem_contents[14'h1ca7] = 8'he4;
s_mem_contents[14'h1ca8] = 8'h0d;
s_mem_contents[14'h1ca9] = 8'h08;
s_mem_contents[14'h1caa] = 8'h68;
s_mem_contents[14'h1cab] = 8'h48;
s_mem_contents[14'h1cac] = 8'hc9;
s_mem_contents[14'h1cad] = 8'h7d;
s_mem_contents[14'h1cae] = 8'hd0;
s_mem_contents[14'h1caf] = 8'hfe;
s_mem_contents[14'h1cb0] = 8'h28;
s_mem_contents[14'h1cb1] = 8'hca;
s_mem_contents[14'h1cb2] = 8'he4;
s_mem_contents[14'h1cb3] = 8'h0d;
s_mem_contents[14'h1cb4] = 8'h08;
s_mem_contents[14'h1cb5] = 8'h68;
s_mem_contents[14'h1cb6] = 8'h48;
s_mem_contents[14'h1cb7] = 8'hc9;
s_mem_contents[14'h1cb8] = 8'h7f;
s_mem_contents[14'h1cb9] = 8'hd0;
s_mem_contents[14'h1cba] = 8'hfe;
s_mem_contents[14'h1cbb] = 8'h28;
s_mem_contents[14'h1cbc] = 8'hca;
s_mem_contents[14'h1cbd] = 8'he4;
s_mem_contents[14'h1cbe] = 8'h0d;
s_mem_contents[14'h1cbf] = 8'h08;
s_mem_contents[14'h1cc0] = 8'he0;
s_mem_contents[14'h1cc1] = 8'h7e;
s_mem_contents[14'h1cc2] = 8'hd0;
s_mem_contents[14'h1cc3] = 8'hfe;
s_mem_contents[14'h1cc4] = 8'h68;
s_mem_contents[14'h1cc5] = 8'h48;
s_mem_contents[14'h1cc6] = 8'hc9;
s_mem_contents[14'h1cc7] = 8'hfc;
s_mem_contents[14'h1cc8] = 8'hd0;
s_mem_contents[14'h1cc9] = 8'hfe;
s_mem_contents[14'h1cca] = 8'h28;
s_mem_contents[14'h1ccb] = 8'ha9;
s_mem_contents[14'h1ccc] = 8'h00;
s_mem_contents[14'h1ccd] = 8'h48;
s_mem_contents[14'h1cce] = 8'ha2;
s_mem_contents[14'h1ccf] = 8'h80;
s_mem_contents[14'h1cd0] = 8'h28;
s_mem_contents[14'h1cd1] = 8'hec;
s_mem_contents[14'h1cd2] = 8'h1b;
s_mem_contents[14'h1cd3] = 8'h02;
s_mem_contents[14'h1cd4] = 8'h08;
s_mem_contents[14'h1cd5] = 8'h68;
s_mem_contents[14'h1cd6] = 8'h48;
s_mem_contents[14'h1cd7] = 8'hc9;
s_mem_contents[14'h1cd8] = 8'h31;
s_mem_contents[14'h1cd9] = 8'hd0;
s_mem_contents[14'h1cda] = 8'hfe;
s_mem_contents[14'h1cdb] = 8'h28;
s_mem_contents[14'h1cdc] = 8'hca;
s_mem_contents[14'h1cdd] = 8'hec;
s_mem_contents[14'h1cde] = 8'h1b;
s_mem_contents[14'h1cdf] = 8'h02;
s_mem_contents[14'h1ce0] = 8'h08;
s_mem_contents[14'h1ce1] = 8'h68;
s_mem_contents[14'h1ce2] = 8'h48;
s_mem_contents[14'h1ce3] = 8'hc9;
s_mem_contents[14'h1ce4] = 8'h33;
s_mem_contents[14'h1ce5] = 8'hd0;
s_mem_contents[14'h1ce6] = 8'hfe;
s_mem_contents[14'h1ce7] = 8'h28;
s_mem_contents[14'h1ce8] = 8'hca;
s_mem_contents[14'h1ce9] = 8'hec;
s_mem_contents[14'h1cea] = 8'h1b;
s_mem_contents[14'h1ceb] = 8'h02;
s_mem_contents[14'h1cec] = 8'h08;
s_mem_contents[14'h1ced] = 8'he0;
s_mem_contents[14'h1cee] = 8'h7e;
s_mem_contents[14'h1cef] = 8'hd0;
s_mem_contents[14'h1cf0] = 8'hfe;
s_mem_contents[14'h1cf1] = 8'h68;
s_mem_contents[14'h1cf2] = 8'h48;
s_mem_contents[14'h1cf3] = 8'hc9;
s_mem_contents[14'h1cf4] = 8'hb0;
s_mem_contents[14'h1cf5] = 8'hd0;
s_mem_contents[14'h1cf6] = 8'hfe;
s_mem_contents[14'h1cf7] = 8'h28;
s_mem_contents[14'h1cf8] = 8'ha9;
s_mem_contents[14'h1cf9] = 8'hff;
s_mem_contents[14'h1cfa] = 8'h48;
s_mem_contents[14'h1cfb] = 8'ha2;
s_mem_contents[14'h1cfc] = 8'h80;
s_mem_contents[14'h1cfd] = 8'h28;
s_mem_contents[14'h1cfe] = 8'hec;
s_mem_contents[14'h1cff] = 8'h1b;
s_mem_contents[14'h1d00] = 8'h02;
s_mem_contents[14'h1d01] = 8'h08;
s_mem_contents[14'h1d02] = 8'h68;
s_mem_contents[14'h1d03] = 8'h48;
s_mem_contents[14'h1d04] = 8'hc9;
s_mem_contents[14'h1d05] = 8'h7d;
s_mem_contents[14'h1d06] = 8'hd0;
s_mem_contents[14'h1d07] = 8'hfe;
s_mem_contents[14'h1d08] = 8'h28;
s_mem_contents[14'h1d09] = 8'hca;
s_mem_contents[14'h1d0a] = 8'hec;
s_mem_contents[14'h1d0b] = 8'h1b;
s_mem_contents[14'h1d0c] = 8'h02;
s_mem_contents[14'h1d0d] = 8'h08;
s_mem_contents[14'h1d0e] = 8'h68;
s_mem_contents[14'h1d0f] = 8'h48;
s_mem_contents[14'h1d10] = 8'hc9;
s_mem_contents[14'h1d11] = 8'h7f;
s_mem_contents[14'h1d12] = 8'hd0;
s_mem_contents[14'h1d13] = 8'hfe;
s_mem_contents[14'h1d14] = 8'h28;
s_mem_contents[14'h1d15] = 8'hca;
s_mem_contents[14'h1d16] = 8'hec;
s_mem_contents[14'h1d17] = 8'h1b;
s_mem_contents[14'h1d18] = 8'h02;
s_mem_contents[14'h1d19] = 8'h08;
s_mem_contents[14'h1d1a] = 8'he0;
s_mem_contents[14'h1d1b] = 8'h7e;
s_mem_contents[14'h1d1c] = 8'hd0;
s_mem_contents[14'h1d1d] = 8'hfe;
s_mem_contents[14'h1d1e] = 8'h68;
s_mem_contents[14'h1d1f] = 8'h48;
s_mem_contents[14'h1d20] = 8'hc9;
s_mem_contents[14'h1d21] = 8'hfc;
s_mem_contents[14'h1d22] = 8'hd0;
s_mem_contents[14'h1d23] = 8'hfe;
s_mem_contents[14'h1d24] = 8'h28;
s_mem_contents[14'h1d25] = 8'ha9;
s_mem_contents[14'h1d26] = 8'h00;
s_mem_contents[14'h1d27] = 8'h48;
s_mem_contents[14'h1d28] = 8'ha2;
s_mem_contents[14'h1d29] = 8'h80;
s_mem_contents[14'h1d2a] = 8'h28;
s_mem_contents[14'h1d2b] = 8'he0;
s_mem_contents[14'h1d2c] = 8'h7f;
s_mem_contents[14'h1d2d] = 8'h08;
s_mem_contents[14'h1d2e] = 8'h68;
s_mem_contents[14'h1d2f] = 8'h48;
s_mem_contents[14'h1d30] = 8'hc9;
s_mem_contents[14'h1d31] = 8'h31;
s_mem_contents[14'h1d32] = 8'hd0;
s_mem_contents[14'h1d33] = 8'hfe;
s_mem_contents[14'h1d34] = 8'h28;
s_mem_contents[14'h1d35] = 8'hca;
s_mem_contents[14'h1d36] = 8'he0;
s_mem_contents[14'h1d37] = 8'h7f;
s_mem_contents[14'h1d38] = 8'h08;
s_mem_contents[14'h1d39] = 8'h68;
s_mem_contents[14'h1d3a] = 8'h48;
s_mem_contents[14'h1d3b] = 8'hc9;
s_mem_contents[14'h1d3c] = 8'h33;
s_mem_contents[14'h1d3d] = 8'hd0;
s_mem_contents[14'h1d3e] = 8'hfe;
s_mem_contents[14'h1d3f] = 8'h28;
s_mem_contents[14'h1d40] = 8'hca;
s_mem_contents[14'h1d41] = 8'he0;
s_mem_contents[14'h1d42] = 8'h7f;
s_mem_contents[14'h1d43] = 8'h08;
s_mem_contents[14'h1d44] = 8'he0;
s_mem_contents[14'h1d45] = 8'h7e;
s_mem_contents[14'h1d46] = 8'hd0;
s_mem_contents[14'h1d47] = 8'hfe;
s_mem_contents[14'h1d48] = 8'h68;
s_mem_contents[14'h1d49] = 8'h48;
s_mem_contents[14'h1d4a] = 8'hc9;
s_mem_contents[14'h1d4b] = 8'hb0;
s_mem_contents[14'h1d4c] = 8'hd0;
s_mem_contents[14'h1d4d] = 8'hfe;
s_mem_contents[14'h1d4e] = 8'h28;
s_mem_contents[14'h1d4f] = 8'ha9;
s_mem_contents[14'h1d50] = 8'hff;
s_mem_contents[14'h1d51] = 8'h48;
s_mem_contents[14'h1d52] = 8'ha2;
s_mem_contents[14'h1d53] = 8'h80;
s_mem_contents[14'h1d54] = 8'h28;
s_mem_contents[14'h1d55] = 8'he0;
s_mem_contents[14'h1d56] = 8'h7f;
s_mem_contents[14'h1d57] = 8'h08;
s_mem_contents[14'h1d58] = 8'h68;
s_mem_contents[14'h1d59] = 8'h48;
s_mem_contents[14'h1d5a] = 8'hc9;
s_mem_contents[14'h1d5b] = 8'h7d;
s_mem_contents[14'h1d5c] = 8'hd0;
s_mem_contents[14'h1d5d] = 8'hfe;
s_mem_contents[14'h1d5e] = 8'h28;
s_mem_contents[14'h1d5f] = 8'hca;
s_mem_contents[14'h1d60] = 8'he0;
s_mem_contents[14'h1d61] = 8'h7f;
s_mem_contents[14'h1d62] = 8'h08;
s_mem_contents[14'h1d63] = 8'h68;
s_mem_contents[14'h1d64] = 8'h48;
s_mem_contents[14'h1d65] = 8'hc9;
s_mem_contents[14'h1d66] = 8'h7f;
s_mem_contents[14'h1d67] = 8'hd0;
s_mem_contents[14'h1d68] = 8'hfe;
s_mem_contents[14'h1d69] = 8'h28;
s_mem_contents[14'h1d6a] = 8'hca;
s_mem_contents[14'h1d6b] = 8'he0;
s_mem_contents[14'h1d6c] = 8'h7f;
s_mem_contents[14'h1d6d] = 8'h08;
s_mem_contents[14'h1d6e] = 8'he0;
s_mem_contents[14'h1d6f] = 8'h7e;
s_mem_contents[14'h1d70] = 8'hd0;
s_mem_contents[14'h1d71] = 8'hfe;
s_mem_contents[14'h1d72] = 8'h68;
s_mem_contents[14'h1d73] = 8'h48;
s_mem_contents[14'h1d74] = 8'hc9;
s_mem_contents[14'h1d75] = 8'hfc;
s_mem_contents[14'h1d76] = 8'hd0;
s_mem_contents[14'h1d77] = 8'hfe;
s_mem_contents[14'h1d78] = 8'h28;
s_mem_contents[14'h1d79] = 8'had;
s_mem_contents[14'h1d7a] = 8'h00;
s_mem_contents[14'h1d7b] = 8'h02;
s_mem_contents[14'h1d7c] = 8'hc9;
s_mem_contents[14'h1d7d] = 8'h1a;
s_mem_contents[14'h1d7e] = 8'hd0;
s_mem_contents[14'h1d7f] = 8'hfe;
s_mem_contents[14'h1d80] = 8'ha9;
s_mem_contents[14'h1d81] = 8'h1b;
s_mem_contents[14'h1d82] = 8'h8d;
s_mem_contents[14'h1d83] = 8'h00;
s_mem_contents[14'h1d84] = 8'h02;
s_mem_contents[14'h1d85] = 8'ha9;
s_mem_contents[14'h1d86] = 8'h00;
s_mem_contents[14'h1d87] = 8'h48;
s_mem_contents[14'h1d88] = 8'ha0;
s_mem_contents[14'h1d89] = 8'h80;
s_mem_contents[14'h1d8a] = 8'h28;
s_mem_contents[14'h1d8b] = 8'hc4;
s_mem_contents[14'h1d8c] = 8'h0d;
s_mem_contents[14'h1d8d] = 8'h08;
s_mem_contents[14'h1d8e] = 8'h68;
s_mem_contents[14'h1d8f] = 8'h48;
s_mem_contents[14'h1d90] = 8'hc9;
s_mem_contents[14'h1d91] = 8'h31;
s_mem_contents[14'h1d92] = 8'hd0;
s_mem_contents[14'h1d93] = 8'hfe;
s_mem_contents[14'h1d94] = 8'h28;
s_mem_contents[14'h1d95] = 8'h88;
s_mem_contents[14'h1d96] = 8'hc4;
s_mem_contents[14'h1d97] = 8'h0d;
s_mem_contents[14'h1d98] = 8'h08;
s_mem_contents[14'h1d99] = 8'h68;
s_mem_contents[14'h1d9a] = 8'h48;
s_mem_contents[14'h1d9b] = 8'hc9;
s_mem_contents[14'h1d9c] = 8'h33;
s_mem_contents[14'h1d9d] = 8'hd0;
s_mem_contents[14'h1d9e] = 8'hfe;
s_mem_contents[14'h1d9f] = 8'h28;
s_mem_contents[14'h1da0] = 8'h88;
s_mem_contents[14'h1da1] = 8'hc4;
s_mem_contents[14'h1da2] = 8'h0d;
s_mem_contents[14'h1da3] = 8'h08;
s_mem_contents[14'h1da4] = 8'hc0;
s_mem_contents[14'h1da5] = 8'h7e;
s_mem_contents[14'h1da6] = 8'hd0;
s_mem_contents[14'h1da7] = 8'hfe;
s_mem_contents[14'h1da8] = 8'h68;
s_mem_contents[14'h1da9] = 8'h48;
s_mem_contents[14'h1daa] = 8'hc9;
s_mem_contents[14'h1dab] = 8'hb0;
s_mem_contents[14'h1dac] = 8'hd0;
s_mem_contents[14'h1dad] = 8'hfe;
s_mem_contents[14'h1dae] = 8'h28;
s_mem_contents[14'h1daf] = 8'ha9;
s_mem_contents[14'h1db0] = 8'hff;
s_mem_contents[14'h1db1] = 8'h48;
s_mem_contents[14'h1db2] = 8'ha0;
s_mem_contents[14'h1db3] = 8'h80;
s_mem_contents[14'h1db4] = 8'h28;
s_mem_contents[14'h1db5] = 8'hc4;
s_mem_contents[14'h1db6] = 8'h0d;
s_mem_contents[14'h1db7] = 8'h08;
s_mem_contents[14'h1db8] = 8'h68;
s_mem_contents[14'h1db9] = 8'h48;
s_mem_contents[14'h1dba] = 8'hc9;
s_mem_contents[14'h1dbb] = 8'h7d;
s_mem_contents[14'h1dbc] = 8'hd0;
s_mem_contents[14'h1dbd] = 8'hfe;
s_mem_contents[14'h1dbe] = 8'h28;
s_mem_contents[14'h1dbf] = 8'h88;
s_mem_contents[14'h1dc0] = 8'hc4;
s_mem_contents[14'h1dc1] = 8'h0d;
s_mem_contents[14'h1dc2] = 8'h08;
s_mem_contents[14'h1dc3] = 8'h68;
s_mem_contents[14'h1dc4] = 8'h48;
s_mem_contents[14'h1dc5] = 8'hc9;
s_mem_contents[14'h1dc6] = 8'h7f;
s_mem_contents[14'h1dc7] = 8'hd0;
s_mem_contents[14'h1dc8] = 8'hfe;
s_mem_contents[14'h1dc9] = 8'h28;
s_mem_contents[14'h1dca] = 8'h88;
s_mem_contents[14'h1dcb] = 8'hc4;
s_mem_contents[14'h1dcc] = 8'h0d;
s_mem_contents[14'h1dcd] = 8'h08;
s_mem_contents[14'h1dce] = 8'hc0;
s_mem_contents[14'h1dcf] = 8'h7e;
s_mem_contents[14'h1dd0] = 8'hd0;
s_mem_contents[14'h1dd1] = 8'hfe;
s_mem_contents[14'h1dd2] = 8'h68;
s_mem_contents[14'h1dd3] = 8'h48;
s_mem_contents[14'h1dd4] = 8'hc9;
s_mem_contents[14'h1dd5] = 8'hfc;
s_mem_contents[14'h1dd6] = 8'hd0;
s_mem_contents[14'h1dd7] = 8'hfe;
s_mem_contents[14'h1dd8] = 8'h28;
s_mem_contents[14'h1dd9] = 8'ha9;
s_mem_contents[14'h1dda] = 8'h00;
s_mem_contents[14'h1ddb] = 8'h48;
s_mem_contents[14'h1ddc] = 8'ha0;
s_mem_contents[14'h1ddd] = 8'h80;
s_mem_contents[14'h1dde] = 8'h28;
s_mem_contents[14'h1ddf] = 8'hcc;
s_mem_contents[14'h1de0] = 8'h1b;
s_mem_contents[14'h1de1] = 8'h02;
s_mem_contents[14'h1de2] = 8'h08;
s_mem_contents[14'h1de3] = 8'h68;
s_mem_contents[14'h1de4] = 8'h48;
s_mem_contents[14'h1de5] = 8'hc9;
s_mem_contents[14'h1de6] = 8'h31;
s_mem_contents[14'h1de7] = 8'hd0;
s_mem_contents[14'h1de8] = 8'hfe;
s_mem_contents[14'h1de9] = 8'h28;
s_mem_contents[14'h1dea] = 8'h88;
s_mem_contents[14'h1deb] = 8'hcc;
s_mem_contents[14'h1dec] = 8'h1b;
s_mem_contents[14'h1ded] = 8'h02;
s_mem_contents[14'h1dee] = 8'h08;
s_mem_contents[14'h1def] = 8'h68;
s_mem_contents[14'h1df0] = 8'h48;
s_mem_contents[14'h1df1] = 8'hc9;
s_mem_contents[14'h1df2] = 8'h33;
s_mem_contents[14'h1df3] = 8'hd0;
s_mem_contents[14'h1df4] = 8'hfe;
s_mem_contents[14'h1df5] = 8'h28;
s_mem_contents[14'h1df6] = 8'h88;
s_mem_contents[14'h1df7] = 8'hcc;
s_mem_contents[14'h1df8] = 8'h1b;
s_mem_contents[14'h1df9] = 8'h02;
s_mem_contents[14'h1dfa] = 8'h08;
s_mem_contents[14'h1dfb] = 8'hc0;
s_mem_contents[14'h1dfc] = 8'h7e;
s_mem_contents[14'h1dfd] = 8'hd0;
s_mem_contents[14'h1dfe] = 8'hfe;
s_mem_contents[14'h1dff] = 8'h68;
s_mem_contents[14'h1e00] = 8'h48;
s_mem_contents[14'h1e01] = 8'hc9;
s_mem_contents[14'h1e02] = 8'hb0;
s_mem_contents[14'h1e03] = 8'hd0;
s_mem_contents[14'h1e04] = 8'hfe;
s_mem_contents[14'h1e05] = 8'h28;
s_mem_contents[14'h1e06] = 8'ha9;
s_mem_contents[14'h1e07] = 8'hff;
s_mem_contents[14'h1e08] = 8'h48;
s_mem_contents[14'h1e09] = 8'ha0;
s_mem_contents[14'h1e0a] = 8'h80;
s_mem_contents[14'h1e0b] = 8'h28;
s_mem_contents[14'h1e0c] = 8'hcc;
s_mem_contents[14'h1e0d] = 8'h1b;
s_mem_contents[14'h1e0e] = 8'h02;
s_mem_contents[14'h1e0f] = 8'h08;
s_mem_contents[14'h1e10] = 8'h68;
s_mem_contents[14'h1e11] = 8'h48;
s_mem_contents[14'h1e12] = 8'hc9;
s_mem_contents[14'h1e13] = 8'h7d;
s_mem_contents[14'h1e14] = 8'hd0;
s_mem_contents[14'h1e15] = 8'hfe;
s_mem_contents[14'h1e16] = 8'h28;
s_mem_contents[14'h1e17] = 8'h88;
s_mem_contents[14'h1e18] = 8'hcc;
s_mem_contents[14'h1e19] = 8'h1b;
s_mem_contents[14'h1e1a] = 8'h02;
s_mem_contents[14'h1e1b] = 8'h08;
s_mem_contents[14'h1e1c] = 8'h68;
s_mem_contents[14'h1e1d] = 8'h48;
s_mem_contents[14'h1e1e] = 8'hc9;
s_mem_contents[14'h1e1f] = 8'h7f;
s_mem_contents[14'h1e20] = 8'hd0;
s_mem_contents[14'h1e21] = 8'hfe;
s_mem_contents[14'h1e22] = 8'h28;
s_mem_contents[14'h1e23] = 8'h88;
s_mem_contents[14'h1e24] = 8'hcc;
s_mem_contents[14'h1e25] = 8'h1b;
s_mem_contents[14'h1e26] = 8'h02;
s_mem_contents[14'h1e27] = 8'h08;
s_mem_contents[14'h1e28] = 8'hc0;
s_mem_contents[14'h1e29] = 8'h7e;
s_mem_contents[14'h1e2a] = 8'hd0;
s_mem_contents[14'h1e2b] = 8'hfe;
s_mem_contents[14'h1e2c] = 8'h68;
s_mem_contents[14'h1e2d] = 8'h48;
s_mem_contents[14'h1e2e] = 8'hc9;
s_mem_contents[14'h1e2f] = 8'hfc;
s_mem_contents[14'h1e30] = 8'hd0;
s_mem_contents[14'h1e31] = 8'hfe;
s_mem_contents[14'h1e32] = 8'h28;
s_mem_contents[14'h1e33] = 8'ha9;
s_mem_contents[14'h1e34] = 8'h00;
s_mem_contents[14'h1e35] = 8'h48;
s_mem_contents[14'h1e36] = 8'ha0;
s_mem_contents[14'h1e37] = 8'h80;
s_mem_contents[14'h1e38] = 8'h28;
s_mem_contents[14'h1e39] = 8'hc0;
s_mem_contents[14'h1e3a] = 8'h7f;
s_mem_contents[14'h1e3b] = 8'h08;
s_mem_contents[14'h1e3c] = 8'h68;
s_mem_contents[14'h1e3d] = 8'h48;
s_mem_contents[14'h1e3e] = 8'hc9;
s_mem_contents[14'h1e3f] = 8'h31;
s_mem_contents[14'h1e40] = 8'hd0;
s_mem_contents[14'h1e41] = 8'hfe;
s_mem_contents[14'h1e42] = 8'h28;
s_mem_contents[14'h1e43] = 8'h88;
s_mem_contents[14'h1e44] = 8'hc0;
s_mem_contents[14'h1e45] = 8'h7f;
s_mem_contents[14'h1e46] = 8'h08;
s_mem_contents[14'h1e47] = 8'h68;
s_mem_contents[14'h1e48] = 8'h48;
s_mem_contents[14'h1e49] = 8'hc9;
s_mem_contents[14'h1e4a] = 8'h33;
s_mem_contents[14'h1e4b] = 8'hd0;
s_mem_contents[14'h1e4c] = 8'hfe;
s_mem_contents[14'h1e4d] = 8'h28;
s_mem_contents[14'h1e4e] = 8'h88;
s_mem_contents[14'h1e4f] = 8'hc0;
s_mem_contents[14'h1e50] = 8'h7f;
s_mem_contents[14'h1e51] = 8'h08;
s_mem_contents[14'h1e52] = 8'hc0;
s_mem_contents[14'h1e53] = 8'h7e;
s_mem_contents[14'h1e54] = 8'hd0;
s_mem_contents[14'h1e55] = 8'hfe;
s_mem_contents[14'h1e56] = 8'h68;
s_mem_contents[14'h1e57] = 8'h48;
s_mem_contents[14'h1e58] = 8'hc9;
s_mem_contents[14'h1e59] = 8'hb0;
s_mem_contents[14'h1e5a] = 8'hd0;
s_mem_contents[14'h1e5b] = 8'hfe;
s_mem_contents[14'h1e5c] = 8'h28;
s_mem_contents[14'h1e5d] = 8'ha9;
s_mem_contents[14'h1e5e] = 8'hff;
s_mem_contents[14'h1e5f] = 8'h48;
s_mem_contents[14'h1e60] = 8'ha0;
s_mem_contents[14'h1e61] = 8'h80;
s_mem_contents[14'h1e62] = 8'h28;
s_mem_contents[14'h1e63] = 8'hc0;
s_mem_contents[14'h1e64] = 8'h7f;
s_mem_contents[14'h1e65] = 8'h08;
s_mem_contents[14'h1e66] = 8'h68;
s_mem_contents[14'h1e67] = 8'h48;
s_mem_contents[14'h1e68] = 8'hc9;
s_mem_contents[14'h1e69] = 8'h7d;
s_mem_contents[14'h1e6a] = 8'hd0;
s_mem_contents[14'h1e6b] = 8'hfe;
s_mem_contents[14'h1e6c] = 8'h28;
s_mem_contents[14'h1e6d] = 8'h88;
s_mem_contents[14'h1e6e] = 8'hc0;
s_mem_contents[14'h1e6f] = 8'h7f;
s_mem_contents[14'h1e70] = 8'h08;
s_mem_contents[14'h1e71] = 8'h68;
s_mem_contents[14'h1e72] = 8'h48;
s_mem_contents[14'h1e73] = 8'hc9;
s_mem_contents[14'h1e74] = 8'h7f;
s_mem_contents[14'h1e75] = 8'hd0;
s_mem_contents[14'h1e76] = 8'hfe;
s_mem_contents[14'h1e77] = 8'h28;
s_mem_contents[14'h1e78] = 8'h88;
s_mem_contents[14'h1e79] = 8'hc0;
s_mem_contents[14'h1e7a] = 8'h7f;
s_mem_contents[14'h1e7b] = 8'h08;
s_mem_contents[14'h1e7c] = 8'hc0;
s_mem_contents[14'h1e7d] = 8'h7e;
s_mem_contents[14'h1e7e] = 8'hd0;
s_mem_contents[14'h1e7f] = 8'hfe;
s_mem_contents[14'h1e80] = 8'h68;
s_mem_contents[14'h1e81] = 8'h48;
s_mem_contents[14'h1e82] = 8'hc9;
s_mem_contents[14'h1e83] = 8'hfc;
s_mem_contents[14'h1e84] = 8'hd0;
s_mem_contents[14'h1e85] = 8'hfe;
s_mem_contents[14'h1e86] = 8'h28;
s_mem_contents[14'h1e87] = 8'had;
s_mem_contents[14'h1e88] = 8'h00;
s_mem_contents[14'h1e89] = 8'h02;
s_mem_contents[14'h1e8a] = 8'hc9;
s_mem_contents[14'h1e8b] = 8'h1b;
s_mem_contents[14'h1e8c] = 8'hd0;
s_mem_contents[14'h1e8d] = 8'hfe;
s_mem_contents[14'h1e8e] = 8'ha9;
s_mem_contents[14'h1e8f] = 8'h1c;
s_mem_contents[14'h1e90] = 8'h8d;
s_mem_contents[14'h1e91] = 8'h00;
s_mem_contents[14'h1e92] = 8'h02;
s_mem_contents[14'h1e93] = 8'ha9;
s_mem_contents[14'h1e94] = 8'h00;
s_mem_contents[14'h1e95] = 8'h48;
s_mem_contents[14'h1e96] = 8'ha9;
s_mem_contents[14'h1e97] = 8'h80;
s_mem_contents[14'h1e98] = 8'h28;
s_mem_contents[14'h1e99] = 8'hc5;
s_mem_contents[14'h1e9a] = 8'h0d;
s_mem_contents[14'h1e9b] = 8'h08;
s_mem_contents[14'h1e9c] = 8'hc9;
s_mem_contents[14'h1e9d] = 8'h80;
s_mem_contents[14'h1e9e] = 8'hd0;
s_mem_contents[14'h1e9f] = 8'hfe;
s_mem_contents[14'h1ea0] = 8'h68;
s_mem_contents[14'h1ea1] = 8'h48;
s_mem_contents[14'h1ea2] = 8'hc9;
s_mem_contents[14'h1ea3] = 8'h31;
s_mem_contents[14'h1ea4] = 8'hd0;
s_mem_contents[14'h1ea5] = 8'hfe;
s_mem_contents[14'h1ea6] = 8'h28;
s_mem_contents[14'h1ea7] = 8'ha9;
s_mem_contents[14'h1ea8] = 8'h00;
s_mem_contents[14'h1ea9] = 8'h48;
s_mem_contents[14'h1eaa] = 8'ha9;
s_mem_contents[14'h1eab] = 8'h7f;
s_mem_contents[14'h1eac] = 8'h28;
s_mem_contents[14'h1ead] = 8'hc5;
s_mem_contents[14'h1eae] = 8'h0d;
s_mem_contents[14'h1eaf] = 8'h08;
s_mem_contents[14'h1eb0] = 8'hc9;
s_mem_contents[14'h1eb1] = 8'h7f;
s_mem_contents[14'h1eb2] = 8'hd0;
s_mem_contents[14'h1eb3] = 8'hfe;
s_mem_contents[14'h1eb4] = 8'h68;
s_mem_contents[14'h1eb5] = 8'h48;
s_mem_contents[14'h1eb6] = 8'hc9;
s_mem_contents[14'h1eb7] = 8'h33;
s_mem_contents[14'h1eb8] = 8'hd0;
s_mem_contents[14'h1eb9] = 8'hfe;
s_mem_contents[14'h1eba] = 8'h28;
s_mem_contents[14'h1ebb] = 8'ha9;
s_mem_contents[14'h1ebc] = 8'h00;
s_mem_contents[14'h1ebd] = 8'h48;
s_mem_contents[14'h1ebe] = 8'ha9;
s_mem_contents[14'h1ebf] = 8'h7e;
s_mem_contents[14'h1ec0] = 8'h28;
s_mem_contents[14'h1ec1] = 8'hc5;
s_mem_contents[14'h1ec2] = 8'h0d;
s_mem_contents[14'h1ec3] = 8'h08;
s_mem_contents[14'h1ec4] = 8'hc9;
s_mem_contents[14'h1ec5] = 8'h7e;
s_mem_contents[14'h1ec6] = 8'hd0;
s_mem_contents[14'h1ec7] = 8'hfe;
s_mem_contents[14'h1ec8] = 8'h68;
s_mem_contents[14'h1ec9] = 8'h48;
s_mem_contents[14'h1eca] = 8'hc9;
s_mem_contents[14'h1ecb] = 8'hb0;
s_mem_contents[14'h1ecc] = 8'hd0;
s_mem_contents[14'h1ecd] = 8'hfe;
s_mem_contents[14'h1ece] = 8'h28;
s_mem_contents[14'h1ecf] = 8'ha9;
s_mem_contents[14'h1ed0] = 8'hff;
s_mem_contents[14'h1ed1] = 8'h48;
s_mem_contents[14'h1ed2] = 8'ha9;
s_mem_contents[14'h1ed3] = 8'h80;
s_mem_contents[14'h1ed4] = 8'h28;
s_mem_contents[14'h1ed5] = 8'hc5;
s_mem_contents[14'h1ed6] = 8'h0d;
s_mem_contents[14'h1ed7] = 8'h08;
s_mem_contents[14'h1ed8] = 8'hc9;
s_mem_contents[14'h1ed9] = 8'h80;
s_mem_contents[14'h1eda] = 8'hd0;
s_mem_contents[14'h1edb] = 8'hfe;
s_mem_contents[14'h1edc] = 8'h68;
s_mem_contents[14'h1edd] = 8'h48;
s_mem_contents[14'h1ede] = 8'hc9;
s_mem_contents[14'h1edf] = 8'h7d;
s_mem_contents[14'h1ee0] = 8'hd0;
s_mem_contents[14'h1ee1] = 8'hfe;
s_mem_contents[14'h1ee2] = 8'h28;
s_mem_contents[14'h1ee3] = 8'ha9;
s_mem_contents[14'h1ee4] = 8'hff;
s_mem_contents[14'h1ee5] = 8'h48;
s_mem_contents[14'h1ee6] = 8'ha9;
s_mem_contents[14'h1ee7] = 8'h7f;
s_mem_contents[14'h1ee8] = 8'h28;
s_mem_contents[14'h1ee9] = 8'hc5;
s_mem_contents[14'h1eea] = 8'h0d;
s_mem_contents[14'h1eeb] = 8'h08;
s_mem_contents[14'h1eec] = 8'hc9;
s_mem_contents[14'h1eed] = 8'h7f;
s_mem_contents[14'h1eee] = 8'hd0;
s_mem_contents[14'h1eef] = 8'hfe;
s_mem_contents[14'h1ef0] = 8'h68;
s_mem_contents[14'h1ef1] = 8'h48;
s_mem_contents[14'h1ef2] = 8'hc9;
s_mem_contents[14'h1ef3] = 8'h7f;
s_mem_contents[14'h1ef4] = 8'hd0;
s_mem_contents[14'h1ef5] = 8'hfe;
s_mem_contents[14'h1ef6] = 8'h28;
s_mem_contents[14'h1ef7] = 8'ha9;
s_mem_contents[14'h1ef8] = 8'hff;
s_mem_contents[14'h1ef9] = 8'h48;
s_mem_contents[14'h1efa] = 8'ha9;
s_mem_contents[14'h1efb] = 8'h7e;
s_mem_contents[14'h1efc] = 8'h28;
s_mem_contents[14'h1efd] = 8'hc5;
s_mem_contents[14'h1efe] = 8'h0d;
s_mem_contents[14'h1eff] = 8'h08;
s_mem_contents[14'h1f00] = 8'hc9;
s_mem_contents[14'h1f01] = 8'h7e;
s_mem_contents[14'h1f02] = 8'hd0;
s_mem_contents[14'h1f03] = 8'hfe;
s_mem_contents[14'h1f04] = 8'h68;
s_mem_contents[14'h1f05] = 8'h48;
s_mem_contents[14'h1f06] = 8'hc9;
s_mem_contents[14'h1f07] = 8'hfc;
s_mem_contents[14'h1f08] = 8'hd0;
s_mem_contents[14'h1f09] = 8'hfe;
s_mem_contents[14'h1f0a] = 8'h28;
s_mem_contents[14'h1f0b] = 8'ha9;
s_mem_contents[14'h1f0c] = 8'h00;
s_mem_contents[14'h1f0d] = 8'h48;
s_mem_contents[14'h1f0e] = 8'ha9;
s_mem_contents[14'h1f0f] = 8'h80;
s_mem_contents[14'h1f10] = 8'h28;
s_mem_contents[14'h1f11] = 8'hcd;
s_mem_contents[14'h1f12] = 8'h1b;
s_mem_contents[14'h1f13] = 8'h02;
s_mem_contents[14'h1f14] = 8'h08;
s_mem_contents[14'h1f15] = 8'hc9;
s_mem_contents[14'h1f16] = 8'h80;
s_mem_contents[14'h1f17] = 8'hd0;
s_mem_contents[14'h1f18] = 8'hfe;
s_mem_contents[14'h1f19] = 8'h68;
s_mem_contents[14'h1f1a] = 8'h48;
s_mem_contents[14'h1f1b] = 8'hc9;
s_mem_contents[14'h1f1c] = 8'h31;
s_mem_contents[14'h1f1d] = 8'hd0;
s_mem_contents[14'h1f1e] = 8'hfe;
s_mem_contents[14'h1f1f] = 8'h28;
s_mem_contents[14'h1f20] = 8'ha9;
s_mem_contents[14'h1f21] = 8'h00;
s_mem_contents[14'h1f22] = 8'h48;
s_mem_contents[14'h1f23] = 8'ha9;
s_mem_contents[14'h1f24] = 8'h7f;
s_mem_contents[14'h1f25] = 8'h28;
s_mem_contents[14'h1f26] = 8'hcd;
s_mem_contents[14'h1f27] = 8'h1b;
s_mem_contents[14'h1f28] = 8'h02;
s_mem_contents[14'h1f29] = 8'h08;
s_mem_contents[14'h1f2a] = 8'hc9;
s_mem_contents[14'h1f2b] = 8'h7f;
s_mem_contents[14'h1f2c] = 8'hd0;
s_mem_contents[14'h1f2d] = 8'hfe;
s_mem_contents[14'h1f2e] = 8'h68;
s_mem_contents[14'h1f2f] = 8'h48;
s_mem_contents[14'h1f30] = 8'hc9;
s_mem_contents[14'h1f31] = 8'h33;
s_mem_contents[14'h1f32] = 8'hd0;
s_mem_contents[14'h1f33] = 8'hfe;
s_mem_contents[14'h1f34] = 8'h28;
s_mem_contents[14'h1f35] = 8'ha9;
s_mem_contents[14'h1f36] = 8'h00;
s_mem_contents[14'h1f37] = 8'h48;
s_mem_contents[14'h1f38] = 8'ha9;
s_mem_contents[14'h1f39] = 8'h7e;
s_mem_contents[14'h1f3a] = 8'h28;
s_mem_contents[14'h1f3b] = 8'hcd;
s_mem_contents[14'h1f3c] = 8'h1b;
s_mem_contents[14'h1f3d] = 8'h02;
s_mem_contents[14'h1f3e] = 8'h08;
s_mem_contents[14'h1f3f] = 8'hc9;
s_mem_contents[14'h1f40] = 8'h7e;
s_mem_contents[14'h1f41] = 8'hd0;
s_mem_contents[14'h1f42] = 8'hfe;
s_mem_contents[14'h1f43] = 8'h68;
s_mem_contents[14'h1f44] = 8'h48;
s_mem_contents[14'h1f45] = 8'hc9;
s_mem_contents[14'h1f46] = 8'hb0;
s_mem_contents[14'h1f47] = 8'hd0;
s_mem_contents[14'h1f48] = 8'hfe;
s_mem_contents[14'h1f49] = 8'h28;
s_mem_contents[14'h1f4a] = 8'ha9;
s_mem_contents[14'h1f4b] = 8'hff;
s_mem_contents[14'h1f4c] = 8'h48;
s_mem_contents[14'h1f4d] = 8'ha9;
s_mem_contents[14'h1f4e] = 8'h80;
s_mem_contents[14'h1f4f] = 8'h28;
s_mem_contents[14'h1f50] = 8'hcd;
s_mem_contents[14'h1f51] = 8'h1b;
s_mem_contents[14'h1f52] = 8'h02;
s_mem_contents[14'h1f53] = 8'h08;
s_mem_contents[14'h1f54] = 8'hc9;
s_mem_contents[14'h1f55] = 8'h80;
s_mem_contents[14'h1f56] = 8'hd0;
s_mem_contents[14'h1f57] = 8'hfe;
s_mem_contents[14'h1f58] = 8'h68;
s_mem_contents[14'h1f59] = 8'h48;
s_mem_contents[14'h1f5a] = 8'hc9;
s_mem_contents[14'h1f5b] = 8'h7d;
s_mem_contents[14'h1f5c] = 8'hd0;
s_mem_contents[14'h1f5d] = 8'hfe;
s_mem_contents[14'h1f5e] = 8'h28;
s_mem_contents[14'h1f5f] = 8'ha9;
s_mem_contents[14'h1f60] = 8'hff;
s_mem_contents[14'h1f61] = 8'h48;
s_mem_contents[14'h1f62] = 8'ha9;
s_mem_contents[14'h1f63] = 8'h7f;
s_mem_contents[14'h1f64] = 8'h28;
s_mem_contents[14'h1f65] = 8'hcd;
s_mem_contents[14'h1f66] = 8'h1b;
s_mem_contents[14'h1f67] = 8'h02;
s_mem_contents[14'h1f68] = 8'h08;
s_mem_contents[14'h1f69] = 8'hc9;
s_mem_contents[14'h1f6a] = 8'h7f;
s_mem_contents[14'h1f6b] = 8'hd0;
s_mem_contents[14'h1f6c] = 8'hfe;
s_mem_contents[14'h1f6d] = 8'h68;
s_mem_contents[14'h1f6e] = 8'h48;
s_mem_contents[14'h1f6f] = 8'hc9;
s_mem_contents[14'h1f70] = 8'h7f;
s_mem_contents[14'h1f71] = 8'hd0;
s_mem_contents[14'h1f72] = 8'hfe;
s_mem_contents[14'h1f73] = 8'h28;
s_mem_contents[14'h1f74] = 8'ha9;
s_mem_contents[14'h1f75] = 8'hff;
s_mem_contents[14'h1f76] = 8'h48;
s_mem_contents[14'h1f77] = 8'ha9;
s_mem_contents[14'h1f78] = 8'h7e;
s_mem_contents[14'h1f79] = 8'h28;
s_mem_contents[14'h1f7a] = 8'hcd;
s_mem_contents[14'h1f7b] = 8'h1b;
s_mem_contents[14'h1f7c] = 8'h02;
s_mem_contents[14'h1f7d] = 8'h08;
s_mem_contents[14'h1f7e] = 8'hc9;
s_mem_contents[14'h1f7f] = 8'h7e;
s_mem_contents[14'h1f80] = 8'hd0;
s_mem_contents[14'h1f81] = 8'hfe;
s_mem_contents[14'h1f82] = 8'h68;
s_mem_contents[14'h1f83] = 8'h48;
s_mem_contents[14'h1f84] = 8'hc9;
s_mem_contents[14'h1f85] = 8'hfc;
s_mem_contents[14'h1f86] = 8'hd0;
s_mem_contents[14'h1f87] = 8'hfe;
s_mem_contents[14'h1f88] = 8'h28;
s_mem_contents[14'h1f89] = 8'ha9;
s_mem_contents[14'h1f8a] = 8'h00;
s_mem_contents[14'h1f8b] = 8'h48;
s_mem_contents[14'h1f8c] = 8'ha9;
s_mem_contents[14'h1f8d] = 8'h80;
s_mem_contents[14'h1f8e] = 8'h28;
s_mem_contents[14'h1f8f] = 8'hc9;
s_mem_contents[14'h1f90] = 8'h7f;
s_mem_contents[14'h1f91] = 8'h08;
s_mem_contents[14'h1f92] = 8'hc9;
s_mem_contents[14'h1f93] = 8'h80;
s_mem_contents[14'h1f94] = 8'hd0;
s_mem_contents[14'h1f95] = 8'hfe;
s_mem_contents[14'h1f96] = 8'h68;
s_mem_contents[14'h1f97] = 8'h48;
s_mem_contents[14'h1f98] = 8'hc9;
s_mem_contents[14'h1f99] = 8'h31;
s_mem_contents[14'h1f9a] = 8'hd0;
s_mem_contents[14'h1f9b] = 8'hfe;
s_mem_contents[14'h1f9c] = 8'h28;
s_mem_contents[14'h1f9d] = 8'ha9;
s_mem_contents[14'h1f9e] = 8'h00;
s_mem_contents[14'h1f9f] = 8'h48;
s_mem_contents[14'h1fa0] = 8'ha9;
s_mem_contents[14'h1fa1] = 8'h7f;
s_mem_contents[14'h1fa2] = 8'h28;
s_mem_contents[14'h1fa3] = 8'hc9;
s_mem_contents[14'h1fa4] = 8'h7f;
s_mem_contents[14'h1fa5] = 8'h08;
s_mem_contents[14'h1fa6] = 8'hc9;
s_mem_contents[14'h1fa7] = 8'h7f;
s_mem_contents[14'h1fa8] = 8'hd0;
s_mem_contents[14'h1fa9] = 8'hfe;
s_mem_contents[14'h1faa] = 8'h68;
s_mem_contents[14'h1fab] = 8'h48;
s_mem_contents[14'h1fac] = 8'hc9;
s_mem_contents[14'h1fad] = 8'h33;
s_mem_contents[14'h1fae] = 8'hd0;
s_mem_contents[14'h1faf] = 8'hfe;
s_mem_contents[14'h1fb0] = 8'h28;
s_mem_contents[14'h1fb1] = 8'ha9;
s_mem_contents[14'h1fb2] = 8'h00;
s_mem_contents[14'h1fb3] = 8'h48;
s_mem_contents[14'h1fb4] = 8'ha9;
s_mem_contents[14'h1fb5] = 8'h7e;
s_mem_contents[14'h1fb6] = 8'h28;
s_mem_contents[14'h1fb7] = 8'hc9;
s_mem_contents[14'h1fb8] = 8'h7f;
s_mem_contents[14'h1fb9] = 8'h08;
s_mem_contents[14'h1fba] = 8'hc9;
s_mem_contents[14'h1fbb] = 8'h7e;
s_mem_contents[14'h1fbc] = 8'hd0;
s_mem_contents[14'h1fbd] = 8'hfe;
s_mem_contents[14'h1fbe] = 8'h68;
s_mem_contents[14'h1fbf] = 8'h48;
s_mem_contents[14'h1fc0] = 8'hc9;
s_mem_contents[14'h1fc1] = 8'hb0;
s_mem_contents[14'h1fc2] = 8'hd0;
s_mem_contents[14'h1fc3] = 8'hfe;
s_mem_contents[14'h1fc4] = 8'h28;
s_mem_contents[14'h1fc5] = 8'ha9;
s_mem_contents[14'h1fc6] = 8'hff;
s_mem_contents[14'h1fc7] = 8'h48;
s_mem_contents[14'h1fc8] = 8'ha9;
s_mem_contents[14'h1fc9] = 8'h80;
s_mem_contents[14'h1fca] = 8'h28;
s_mem_contents[14'h1fcb] = 8'hc9;
s_mem_contents[14'h1fcc] = 8'h7f;
s_mem_contents[14'h1fcd] = 8'h08;
s_mem_contents[14'h1fce] = 8'hc9;
s_mem_contents[14'h1fcf] = 8'h80;
s_mem_contents[14'h1fd0] = 8'hd0;
s_mem_contents[14'h1fd1] = 8'hfe;
s_mem_contents[14'h1fd2] = 8'h68;
s_mem_contents[14'h1fd3] = 8'h48;
s_mem_contents[14'h1fd4] = 8'hc9;
s_mem_contents[14'h1fd5] = 8'h7d;
s_mem_contents[14'h1fd6] = 8'hd0;
s_mem_contents[14'h1fd7] = 8'hfe;
s_mem_contents[14'h1fd8] = 8'h28;
s_mem_contents[14'h1fd9] = 8'ha9;
s_mem_contents[14'h1fda] = 8'hff;
s_mem_contents[14'h1fdb] = 8'h48;
s_mem_contents[14'h1fdc] = 8'ha9;
s_mem_contents[14'h1fdd] = 8'h7f;
s_mem_contents[14'h1fde] = 8'h28;
s_mem_contents[14'h1fdf] = 8'hc9;
s_mem_contents[14'h1fe0] = 8'h7f;
s_mem_contents[14'h1fe1] = 8'h08;
s_mem_contents[14'h1fe2] = 8'hc9;
s_mem_contents[14'h1fe3] = 8'h7f;
s_mem_contents[14'h1fe4] = 8'hd0;
s_mem_contents[14'h1fe5] = 8'hfe;
s_mem_contents[14'h1fe6] = 8'h68;
s_mem_contents[14'h1fe7] = 8'h48;
s_mem_contents[14'h1fe8] = 8'hc9;
s_mem_contents[14'h1fe9] = 8'h7f;
s_mem_contents[14'h1fea] = 8'hd0;
s_mem_contents[14'h1feb] = 8'hfe;
s_mem_contents[14'h1fec] = 8'h28;
s_mem_contents[14'h1fed] = 8'ha9;
s_mem_contents[14'h1fee] = 8'hff;
s_mem_contents[14'h1fef] = 8'h48;
s_mem_contents[14'h1ff0] = 8'ha9;
s_mem_contents[14'h1ff1] = 8'h7e;
s_mem_contents[14'h1ff2] = 8'h28;
s_mem_contents[14'h1ff3] = 8'hc9;
s_mem_contents[14'h1ff4] = 8'h7f;
s_mem_contents[14'h1ff5] = 8'h08;
s_mem_contents[14'h1ff6] = 8'hc9;
s_mem_contents[14'h1ff7] = 8'h7e;
s_mem_contents[14'h1ff8] = 8'hd0;
s_mem_contents[14'h1ff9] = 8'hfe;
s_mem_contents[14'h1ffa] = 8'h68;
s_mem_contents[14'h1ffb] = 8'h48;
s_mem_contents[14'h1ffc] = 8'hc9;
s_mem_contents[14'h1ffd] = 8'hfc;
s_mem_contents[14'h1ffe] = 8'hd0;
s_mem_contents[14'h1fff] = 8'hfe;
s_mem_contents[14'h2000] = 8'h28;
s_mem_contents[14'h2001] = 8'ha2;
s_mem_contents[14'h2002] = 8'h04;
s_mem_contents[14'h2003] = 8'ha9;
s_mem_contents[14'h2004] = 8'h00;
s_mem_contents[14'h2005] = 8'h48;
s_mem_contents[14'h2006] = 8'ha9;
s_mem_contents[14'h2007] = 8'h80;
s_mem_contents[14'h2008] = 8'h28;
s_mem_contents[14'h2009] = 8'hd5;
s_mem_contents[14'h200a] = 8'h09;
s_mem_contents[14'h200b] = 8'h08;
s_mem_contents[14'h200c] = 8'hc9;
s_mem_contents[14'h200d] = 8'h80;
s_mem_contents[14'h200e] = 8'hd0;
s_mem_contents[14'h200f] = 8'hfe;
s_mem_contents[14'h2010] = 8'h68;
s_mem_contents[14'h2011] = 8'h48;
s_mem_contents[14'h2012] = 8'hc9;
s_mem_contents[14'h2013] = 8'h31;
s_mem_contents[14'h2014] = 8'hd0;
s_mem_contents[14'h2015] = 8'hfe;
s_mem_contents[14'h2016] = 8'h28;
s_mem_contents[14'h2017] = 8'ha9;
s_mem_contents[14'h2018] = 8'h00;
s_mem_contents[14'h2019] = 8'h48;
s_mem_contents[14'h201a] = 8'ha9;
s_mem_contents[14'h201b] = 8'h7f;
s_mem_contents[14'h201c] = 8'h28;
s_mem_contents[14'h201d] = 8'hd5;
s_mem_contents[14'h201e] = 8'h09;
s_mem_contents[14'h201f] = 8'h08;
s_mem_contents[14'h2020] = 8'hc9;
s_mem_contents[14'h2021] = 8'h7f;
s_mem_contents[14'h2022] = 8'hd0;
s_mem_contents[14'h2023] = 8'hfe;
s_mem_contents[14'h2024] = 8'h68;
s_mem_contents[14'h2025] = 8'h48;
s_mem_contents[14'h2026] = 8'hc9;
s_mem_contents[14'h2027] = 8'h33;
s_mem_contents[14'h2028] = 8'hd0;
s_mem_contents[14'h2029] = 8'hfe;
s_mem_contents[14'h202a] = 8'h28;
s_mem_contents[14'h202b] = 8'ha9;
s_mem_contents[14'h202c] = 8'h00;
s_mem_contents[14'h202d] = 8'h48;
s_mem_contents[14'h202e] = 8'ha9;
s_mem_contents[14'h202f] = 8'h7e;
s_mem_contents[14'h2030] = 8'h28;
s_mem_contents[14'h2031] = 8'hd5;
s_mem_contents[14'h2032] = 8'h09;
s_mem_contents[14'h2033] = 8'h08;
s_mem_contents[14'h2034] = 8'hc9;
s_mem_contents[14'h2035] = 8'h7e;
s_mem_contents[14'h2036] = 8'hd0;
s_mem_contents[14'h2037] = 8'hfe;
s_mem_contents[14'h2038] = 8'h68;
s_mem_contents[14'h2039] = 8'h48;
s_mem_contents[14'h203a] = 8'hc9;
s_mem_contents[14'h203b] = 8'hb0;
s_mem_contents[14'h203c] = 8'hd0;
s_mem_contents[14'h203d] = 8'hfe;
s_mem_contents[14'h203e] = 8'h28;
s_mem_contents[14'h203f] = 8'ha9;
s_mem_contents[14'h2040] = 8'hff;
s_mem_contents[14'h2041] = 8'h48;
s_mem_contents[14'h2042] = 8'ha9;
s_mem_contents[14'h2043] = 8'h80;
s_mem_contents[14'h2044] = 8'h28;
s_mem_contents[14'h2045] = 8'hd5;
s_mem_contents[14'h2046] = 8'h09;
s_mem_contents[14'h2047] = 8'h08;
s_mem_contents[14'h2048] = 8'hc9;
s_mem_contents[14'h2049] = 8'h80;
s_mem_contents[14'h204a] = 8'hd0;
s_mem_contents[14'h204b] = 8'hfe;
s_mem_contents[14'h204c] = 8'h68;
s_mem_contents[14'h204d] = 8'h48;
s_mem_contents[14'h204e] = 8'hc9;
s_mem_contents[14'h204f] = 8'h7d;
s_mem_contents[14'h2050] = 8'hd0;
s_mem_contents[14'h2051] = 8'hfe;
s_mem_contents[14'h2052] = 8'h28;
s_mem_contents[14'h2053] = 8'ha9;
s_mem_contents[14'h2054] = 8'hff;
s_mem_contents[14'h2055] = 8'h48;
s_mem_contents[14'h2056] = 8'ha9;
s_mem_contents[14'h2057] = 8'h7f;
s_mem_contents[14'h2058] = 8'h28;
s_mem_contents[14'h2059] = 8'hd5;
s_mem_contents[14'h205a] = 8'h09;
s_mem_contents[14'h205b] = 8'h08;
s_mem_contents[14'h205c] = 8'hc9;
s_mem_contents[14'h205d] = 8'h7f;
s_mem_contents[14'h205e] = 8'hd0;
s_mem_contents[14'h205f] = 8'hfe;
s_mem_contents[14'h2060] = 8'h68;
s_mem_contents[14'h2061] = 8'h48;
s_mem_contents[14'h2062] = 8'hc9;
s_mem_contents[14'h2063] = 8'h7f;
s_mem_contents[14'h2064] = 8'hd0;
s_mem_contents[14'h2065] = 8'hfe;
s_mem_contents[14'h2066] = 8'h28;
s_mem_contents[14'h2067] = 8'ha9;
s_mem_contents[14'h2068] = 8'hff;
s_mem_contents[14'h2069] = 8'h48;
s_mem_contents[14'h206a] = 8'ha9;
s_mem_contents[14'h206b] = 8'h7e;
s_mem_contents[14'h206c] = 8'h28;
s_mem_contents[14'h206d] = 8'hd5;
s_mem_contents[14'h206e] = 8'h09;
s_mem_contents[14'h206f] = 8'h08;
s_mem_contents[14'h2070] = 8'hc9;
s_mem_contents[14'h2071] = 8'h7e;
s_mem_contents[14'h2072] = 8'hd0;
s_mem_contents[14'h2073] = 8'hfe;
s_mem_contents[14'h2074] = 8'h68;
s_mem_contents[14'h2075] = 8'h48;
s_mem_contents[14'h2076] = 8'hc9;
s_mem_contents[14'h2077] = 8'hfc;
s_mem_contents[14'h2078] = 8'hd0;
s_mem_contents[14'h2079] = 8'hfe;
s_mem_contents[14'h207a] = 8'h28;
s_mem_contents[14'h207b] = 8'ha9;
s_mem_contents[14'h207c] = 8'h00;
s_mem_contents[14'h207d] = 8'h48;
s_mem_contents[14'h207e] = 8'ha9;
s_mem_contents[14'h207f] = 8'h80;
s_mem_contents[14'h2080] = 8'h28;
s_mem_contents[14'h2081] = 8'hdd;
s_mem_contents[14'h2082] = 8'h17;
s_mem_contents[14'h2083] = 8'h02;
s_mem_contents[14'h2084] = 8'h08;
s_mem_contents[14'h2085] = 8'hc9;
s_mem_contents[14'h2086] = 8'h80;
s_mem_contents[14'h2087] = 8'hd0;
s_mem_contents[14'h2088] = 8'hfe;
s_mem_contents[14'h2089] = 8'h68;
s_mem_contents[14'h208a] = 8'h48;
s_mem_contents[14'h208b] = 8'hc9;
s_mem_contents[14'h208c] = 8'h31;
s_mem_contents[14'h208d] = 8'hd0;
s_mem_contents[14'h208e] = 8'hfe;
s_mem_contents[14'h208f] = 8'h28;
s_mem_contents[14'h2090] = 8'ha9;
s_mem_contents[14'h2091] = 8'h00;
s_mem_contents[14'h2092] = 8'h48;
s_mem_contents[14'h2093] = 8'ha9;
s_mem_contents[14'h2094] = 8'h7f;
s_mem_contents[14'h2095] = 8'h28;
s_mem_contents[14'h2096] = 8'hdd;
s_mem_contents[14'h2097] = 8'h17;
s_mem_contents[14'h2098] = 8'h02;
s_mem_contents[14'h2099] = 8'h08;
s_mem_contents[14'h209a] = 8'hc9;
s_mem_contents[14'h209b] = 8'h7f;
s_mem_contents[14'h209c] = 8'hd0;
s_mem_contents[14'h209d] = 8'hfe;
s_mem_contents[14'h209e] = 8'h68;
s_mem_contents[14'h209f] = 8'h48;
s_mem_contents[14'h20a0] = 8'hc9;
s_mem_contents[14'h20a1] = 8'h33;
s_mem_contents[14'h20a2] = 8'hd0;
s_mem_contents[14'h20a3] = 8'hfe;
s_mem_contents[14'h20a4] = 8'h28;
s_mem_contents[14'h20a5] = 8'ha9;
s_mem_contents[14'h20a6] = 8'h00;
s_mem_contents[14'h20a7] = 8'h48;
s_mem_contents[14'h20a8] = 8'ha9;
s_mem_contents[14'h20a9] = 8'h7e;
s_mem_contents[14'h20aa] = 8'h28;
s_mem_contents[14'h20ab] = 8'hdd;
s_mem_contents[14'h20ac] = 8'h17;
s_mem_contents[14'h20ad] = 8'h02;
s_mem_contents[14'h20ae] = 8'h08;
s_mem_contents[14'h20af] = 8'hc9;
s_mem_contents[14'h20b0] = 8'h7e;
s_mem_contents[14'h20b1] = 8'hd0;
s_mem_contents[14'h20b2] = 8'hfe;
s_mem_contents[14'h20b3] = 8'h68;
s_mem_contents[14'h20b4] = 8'h48;
s_mem_contents[14'h20b5] = 8'hc9;
s_mem_contents[14'h20b6] = 8'hb0;
s_mem_contents[14'h20b7] = 8'hd0;
s_mem_contents[14'h20b8] = 8'hfe;
s_mem_contents[14'h20b9] = 8'h28;
s_mem_contents[14'h20ba] = 8'ha9;
s_mem_contents[14'h20bb] = 8'hff;
s_mem_contents[14'h20bc] = 8'h48;
s_mem_contents[14'h20bd] = 8'ha9;
s_mem_contents[14'h20be] = 8'h80;
s_mem_contents[14'h20bf] = 8'h28;
s_mem_contents[14'h20c0] = 8'hdd;
s_mem_contents[14'h20c1] = 8'h17;
s_mem_contents[14'h20c2] = 8'h02;
s_mem_contents[14'h20c3] = 8'h08;
s_mem_contents[14'h20c4] = 8'hc9;
s_mem_contents[14'h20c5] = 8'h80;
s_mem_contents[14'h20c6] = 8'hd0;
s_mem_contents[14'h20c7] = 8'hfe;
s_mem_contents[14'h20c8] = 8'h68;
s_mem_contents[14'h20c9] = 8'h48;
s_mem_contents[14'h20ca] = 8'hc9;
s_mem_contents[14'h20cb] = 8'h7d;
s_mem_contents[14'h20cc] = 8'hd0;
s_mem_contents[14'h20cd] = 8'hfe;
s_mem_contents[14'h20ce] = 8'h28;
s_mem_contents[14'h20cf] = 8'ha9;
s_mem_contents[14'h20d0] = 8'hff;
s_mem_contents[14'h20d1] = 8'h48;
s_mem_contents[14'h20d2] = 8'ha9;
s_mem_contents[14'h20d3] = 8'h7f;
s_mem_contents[14'h20d4] = 8'h28;
s_mem_contents[14'h20d5] = 8'hdd;
s_mem_contents[14'h20d6] = 8'h17;
s_mem_contents[14'h20d7] = 8'h02;
s_mem_contents[14'h20d8] = 8'h08;
s_mem_contents[14'h20d9] = 8'hc9;
s_mem_contents[14'h20da] = 8'h7f;
s_mem_contents[14'h20db] = 8'hd0;
s_mem_contents[14'h20dc] = 8'hfe;
s_mem_contents[14'h20dd] = 8'h68;
s_mem_contents[14'h20de] = 8'h48;
s_mem_contents[14'h20df] = 8'hc9;
s_mem_contents[14'h20e0] = 8'h7f;
s_mem_contents[14'h20e1] = 8'hd0;
s_mem_contents[14'h20e2] = 8'hfe;
s_mem_contents[14'h20e3] = 8'h28;
s_mem_contents[14'h20e4] = 8'ha9;
s_mem_contents[14'h20e5] = 8'hff;
s_mem_contents[14'h20e6] = 8'h48;
s_mem_contents[14'h20e7] = 8'ha9;
s_mem_contents[14'h20e8] = 8'h7e;
s_mem_contents[14'h20e9] = 8'h28;
s_mem_contents[14'h20ea] = 8'hdd;
s_mem_contents[14'h20eb] = 8'h17;
s_mem_contents[14'h20ec] = 8'h02;
s_mem_contents[14'h20ed] = 8'h08;
s_mem_contents[14'h20ee] = 8'hc9;
s_mem_contents[14'h20ef] = 8'h7e;
s_mem_contents[14'h20f0] = 8'hd0;
s_mem_contents[14'h20f1] = 8'hfe;
s_mem_contents[14'h20f2] = 8'h68;
s_mem_contents[14'h20f3] = 8'h48;
s_mem_contents[14'h20f4] = 8'hc9;
s_mem_contents[14'h20f5] = 8'hfc;
s_mem_contents[14'h20f6] = 8'hd0;
s_mem_contents[14'h20f7] = 8'hfe;
s_mem_contents[14'h20f8] = 8'h28;
s_mem_contents[14'h20f9] = 8'ha0;
s_mem_contents[14'h20fa] = 8'h04;
s_mem_contents[14'h20fb] = 8'ha2;
s_mem_contents[14'h20fc] = 8'h08;
s_mem_contents[14'h20fd] = 8'ha9;
s_mem_contents[14'h20fe] = 8'h00;
s_mem_contents[14'h20ff] = 8'h48;
s_mem_contents[14'h2100] = 8'ha9;
s_mem_contents[14'h2101] = 8'h80;
s_mem_contents[14'h2102] = 8'h28;
s_mem_contents[14'h2103] = 8'hd9;
s_mem_contents[14'h2104] = 8'h17;
s_mem_contents[14'h2105] = 8'h02;
s_mem_contents[14'h2106] = 8'h08;
s_mem_contents[14'h2107] = 8'hc9;
s_mem_contents[14'h2108] = 8'h80;
s_mem_contents[14'h2109] = 8'hd0;
s_mem_contents[14'h210a] = 8'hfe;
s_mem_contents[14'h210b] = 8'h68;
s_mem_contents[14'h210c] = 8'h48;
s_mem_contents[14'h210d] = 8'hc9;
s_mem_contents[14'h210e] = 8'h31;
s_mem_contents[14'h210f] = 8'hd0;
s_mem_contents[14'h2110] = 8'hfe;
s_mem_contents[14'h2111] = 8'h28;
s_mem_contents[14'h2112] = 8'ha9;
s_mem_contents[14'h2113] = 8'h00;
s_mem_contents[14'h2114] = 8'h48;
s_mem_contents[14'h2115] = 8'ha9;
s_mem_contents[14'h2116] = 8'h7f;
s_mem_contents[14'h2117] = 8'h28;
s_mem_contents[14'h2118] = 8'hd9;
s_mem_contents[14'h2119] = 8'h17;
s_mem_contents[14'h211a] = 8'h02;
s_mem_contents[14'h211b] = 8'h08;
s_mem_contents[14'h211c] = 8'hc9;
s_mem_contents[14'h211d] = 8'h7f;
s_mem_contents[14'h211e] = 8'hd0;
s_mem_contents[14'h211f] = 8'hfe;
s_mem_contents[14'h2120] = 8'h68;
s_mem_contents[14'h2121] = 8'h48;
s_mem_contents[14'h2122] = 8'hc9;
s_mem_contents[14'h2123] = 8'h33;
s_mem_contents[14'h2124] = 8'hd0;
s_mem_contents[14'h2125] = 8'hfe;
s_mem_contents[14'h2126] = 8'h28;
s_mem_contents[14'h2127] = 8'ha9;
s_mem_contents[14'h2128] = 8'h00;
s_mem_contents[14'h2129] = 8'h48;
s_mem_contents[14'h212a] = 8'ha9;
s_mem_contents[14'h212b] = 8'h7e;
s_mem_contents[14'h212c] = 8'h28;
s_mem_contents[14'h212d] = 8'hd9;
s_mem_contents[14'h212e] = 8'h17;
s_mem_contents[14'h212f] = 8'h02;
s_mem_contents[14'h2130] = 8'h08;
s_mem_contents[14'h2131] = 8'hc9;
s_mem_contents[14'h2132] = 8'h7e;
s_mem_contents[14'h2133] = 8'hd0;
s_mem_contents[14'h2134] = 8'hfe;
s_mem_contents[14'h2135] = 8'h68;
s_mem_contents[14'h2136] = 8'h48;
s_mem_contents[14'h2137] = 8'hc9;
s_mem_contents[14'h2138] = 8'hb0;
s_mem_contents[14'h2139] = 8'hd0;
s_mem_contents[14'h213a] = 8'hfe;
s_mem_contents[14'h213b] = 8'h28;
s_mem_contents[14'h213c] = 8'ha9;
s_mem_contents[14'h213d] = 8'hff;
s_mem_contents[14'h213e] = 8'h48;
s_mem_contents[14'h213f] = 8'ha9;
s_mem_contents[14'h2140] = 8'h80;
s_mem_contents[14'h2141] = 8'h28;
s_mem_contents[14'h2142] = 8'hd9;
s_mem_contents[14'h2143] = 8'h17;
s_mem_contents[14'h2144] = 8'h02;
s_mem_contents[14'h2145] = 8'h08;
s_mem_contents[14'h2146] = 8'hc9;
s_mem_contents[14'h2147] = 8'h80;
s_mem_contents[14'h2148] = 8'hd0;
s_mem_contents[14'h2149] = 8'hfe;
s_mem_contents[14'h214a] = 8'h68;
s_mem_contents[14'h214b] = 8'h48;
s_mem_contents[14'h214c] = 8'hc9;
s_mem_contents[14'h214d] = 8'h7d;
s_mem_contents[14'h214e] = 8'hd0;
s_mem_contents[14'h214f] = 8'hfe;
s_mem_contents[14'h2150] = 8'h28;
s_mem_contents[14'h2151] = 8'ha9;
s_mem_contents[14'h2152] = 8'hff;
s_mem_contents[14'h2153] = 8'h48;
s_mem_contents[14'h2154] = 8'ha9;
s_mem_contents[14'h2155] = 8'h7f;
s_mem_contents[14'h2156] = 8'h28;
s_mem_contents[14'h2157] = 8'hd9;
s_mem_contents[14'h2158] = 8'h17;
s_mem_contents[14'h2159] = 8'h02;
s_mem_contents[14'h215a] = 8'h08;
s_mem_contents[14'h215b] = 8'hc9;
s_mem_contents[14'h215c] = 8'h7f;
s_mem_contents[14'h215d] = 8'hd0;
s_mem_contents[14'h215e] = 8'hfe;
s_mem_contents[14'h215f] = 8'h68;
s_mem_contents[14'h2160] = 8'h48;
s_mem_contents[14'h2161] = 8'hc9;
s_mem_contents[14'h2162] = 8'h7f;
s_mem_contents[14'h2163] = 8'hd0;
s_mem_contents[14'h2164] = 8'hfe;
s_mem_contents[14'h2165] = 8'h28;
s_mem_contents[14'h2166] = 8'ha9;
s_mem_contents[14'h2167] = 8'hff;
s_mem_contents[14'h2168] = 8'h48;
s_mem_contents[14'h2169] = 8'ha9;
s_mem_contents[14'h216a] = 8'h7e;
s_mem_contents[14'h216b] = 8'h28;
s_mem_contents[14'h216c] = 8'hd9;
s_mem_contents[14'h216d] = 8'h17;
s_mem_contents[14'h216e] = 8'h02;
s_mem_contents[14'h216f] = 8'h08;
s_mem_contents[14'h2170] = 8'hc9;
s_mem_contents[14'h2171] = 8'h7e;
s_mem_contents[14'h2172] = 8'hd0;
s_mem_contents[14'h2173] = 8'hfe;
s_mem_contents[14'h2174] = 8'h68;
s_mem_contents[14'h2175] = 8'h48;
s_mem_contents[14'h2176] = 8'hc9;
s_mem_contents[14'h2177] = 8'hfc;
s_mem_contents[14'h2178] = 8'hd0;
s_mem_contents[14'h2179] = 8'hfe;
s_mem_contents[14'h217a] = 8'h28;
s_mem_contents[14'h217b] = 8'ha9;
s_mem_contents[14'h217c] = 8'h00;
s_mem_contents[14'h217d] = 8'h48;
s_mem_contents[14'h217e] = 8'ha9;
s_mem_contents[14'h217f] = 8'h80;
s_mem_contents[14'h2180] = 8'h28;
s_mem_contents[14'h2181] = 8'hc1;
s_mem_contents[14'h2182] = 8'h1a;
s_mem_contents[14'h2183] = 8'h08;
s_mem_contents[14'h2184] = 8'hc9;
s_mem_contents[14'h2185] = 8'h80;
s_mem_contents[14'h2186] = 8'hd0;
s_mem_contents[14'h2187] = 8'hfe;
s_mem_contents[14'h2188] = 8'h68;
s_mem_contents[14'h2189] = 8'h48;
s_mem_contents[14'h218a] = 8'hc9;
s_mem_contents[14'h218b] = 8'h31;
s_mem_contents[14'h218c] = 8'hd0;
s_mem_contents[14'h218d] = 8'hfe;
s_mem_contents[14'h218e] = 8'h28;
s_mem_contents[14'h218f] = 8'ha9;
s_mem_contents[14'h2190] = 8'h00;
s_mem_contents[14'h2191] = 8'h48;
s_mem_contents[14'h2192] = 8'ha9;
s_mem_contents[14'h2193] = 8'h7f;
s_mem_contents[14'h2194] = 8'h28;
s_mem_contents[14'h2195] = 8'hc1;
s_mem_contents[14'h2196] = 8'h1a;
s_mem_contents[14'h2197] = 8'h08;
s_mem_contents[14'h2198] = 8'hc9;
s_mem_contents[14'h2199] = 8'h7f;
s_mem_contents[14'h219a] = 8'hd0;
s_mem_contents[14'h219b] = 8'hfe;
s_mem_contents[14'h219c] = 8'h68;
s_mem_contents[14'h219d] = 8'h48;
s_mem_contents[14'h219e] = 8'hc9;
s_mem_contents[14'h219f] = 8'h33;
s_mem_contents[14'h21a0] = 8'hd0;
s_mem_contents[14'h21a1] = 8'hfe;
s_mem_contents[14'h21a2] = 8'h28;
s_mem_contents[14'h21a3] = 8'ha9;
s_mem_contents[14'h21a4] = 8'h00;
s_mem_contents[14'h21a5] = 8'h48;
s_mem_contents[14'h21a6] = 8'ha9;
s_mem_contents[14'h21a7] = 8'h7e;
s_mem_contents[14'h21a8] = 8'h28;
s_mem_contents[14'h21a9] = 8'hc1;
s_mem_contents[14'h21aa] = 8'h1a;
s_mem_contents[14'h21ab] = 8'h08;
s_mem_contents[14'h21ac] = 8'hc9;
s_mem_contents[14'h21ad] = 8'h7e;
s_mem_contents[14'h21ae] = 8'hd0;
s_mem_contents[14'h21af] = 8'hfe;
s_mem_contents[14'h21b0] = 8'h68;
s_mem_contents[14'h21b1] = 8'h48;
s_mem_contents[14'h21b2] = 8'hc9;
s_mem_contents[14'h21b3] = 8'hb0;
s_mem_contents[14'h21b4] = 8'hd0;
s_mem_contents[14'h21b5] = 8'hfe;
s_mem_contents[14'h21b6] = 8'h28;
s_mem_contents[14'h21b7] = 8'ha9;
s_mem_contents[14'h21b8] = 8'hff;
s_mem_contents[14'h21b9] = 8'h48;
s_mem_contents[14'h21ba] = 8'ha9;
s_mem_contents[14'h21bb] = 8'h80;
s_mem_contents[14'h21bc] = 8'h28;
s_mem_contents[14'h21bd] = 8'hc1;
s_mem_contents[14'h21be] = 8'h1a;
s_mem_contents[14'h21bf] = 8'h08;
s_mem_contents[14'h21c0] = 8'hc9;
s_mem_contents[14'h21c1] = 8'h80;
s_mem_contents[14'h21c2] = 8'hd0;
s_mem_contents[14'h21c3] = 8'hfe;
s_mem_contents[14'h21c4] = 8'h68;
s_mem_contents[14'h21c5] = 8'h48;
s_mem_contents[14'h21c6] = 8'hc9;
s_mem_contents[14'h21c7] = 8'h7d;
s_mem_contents[14'h21c8] = 8'hd0;
s_mem_contents[14'h21c9] = 8'hfe;
s_mem_contents[14'h21ca] = 8'h28;
s_mem_contents[14'h21cb] = 8'ha9;
s_mem_contents[14'h21cc] = 8'hff;
s_mem_contents[14'h21cd] = 8'h48;
s_mem_contents[14'h21ce] = 8'ha9;
s_mem_contents[14'h21cf] = 8'h7f;
s_mem_contents[14'h21d0] = 8'h28;
s_mem_contents[14'h21d1] = 8'hc1;
s_mem_contents[14'h21d2] = 8'h1a;
s_mem_contents[14'h21d3] = 8'h08;
s_mem_contents[14'h21d4] = 8'hc9;
s_mem_contents[14'h21d5] = 8'h7f;
s_mem_contents[14'h21d6] = 8'hd0;
s_mem_contents[14'h21d7] = 8'hfe;
s_mem_contents[14'h21d8] = 8'h68;
s_mem_contents[14'h21d9] = 8'h48;
s_mem_contents[14'h21da] = 8'hc9;
s_mem_contents[14'h21db] = 8'h7f;
s_mem_contents[14'h21dc] = 8'hd0;
s_mem_contents[14'h21dd] = 8'hfe;
s_mem_contents[14'h21de] = 8'h28;
s_mem_contents[14'h21df] = 8'ha9;
s_mem_contents[14'h21e0] = 8'hff;
s_mem_contents[14'h21e1] = 8'h48;
s_mem_contents[14'h21e2] = 8'ha9;
s_mem_contents[14'h21e3] = 8'h7e;
s_mem_contents[14'h21e4] = 8'h28;
s_mem_contents[14'h21e5] = 8'hc1;
s_mem_contents[14'h21e6] = 8'h1a;
s_mem_contents[14'h21e7] = 8'h08;
s_mem_contents[14'h21e8] = 8'hc9;
s_mem_contents[14'h21e9] = 8'h7e;
s_mem_contents[14'h21ea] = 8'hd0;
s_mem_contents[14'h21eb] = 8'hfe;
s_mem_contents[14'h21ec] = 8'h68;
s_mem_contents[14'h21ed] = 8'h48;
s_mem_contents[14'h21ee] = 8'hc9;
s_mem_contents[14'h21ef] = 8'hfc;
s_mem_contents[14'h21f0] = 8'hd0;
s_mem_contents[14'h21f1] = 8'hfe;
s_mem_contents[14'h21f2] = 8'h28;
s_mem_contents[14'h21f3] = 8'ha9;
s_mem_contents[14'h21f4] = 8'h00;
s_mem_contents[14'h21f5] = 8'h48;
s_mem_contents[14'h21f6] = 8'ha9;
s_mem_contents[14'h21f7] = 8'h80;
s_mem_contents[14'h21f8] = 8'h28;
s_mem_contents[14'h21f9] = 8'hd1;
s_mem_contents[14'h21fa] = 8'h1a;
s_mem_contents[14'h21fb] = 8'h08;
s_mem_contents[14'h21fc] = 8'hc9;
s_mem_contents[14'h21fd] = 8'h80;
s_mem_contents[14'h21fe] = 8'hd0;
s_mem_contents[14'h21ff] = 8'hfe;
s_mem_contents[14'h2200] = 8'h68;
s_mem_contents[14'h2201] = 8'h48;
s_mem_contents[14'h2202] = 8'hc9;
s_mem_contents[14'h2203] = 8'h31;
s_mem_contents[14'h2204] = 8'hd0;
s_mem_contents[14'h2205] = 8'hfe;
s_mem_contents[14'h2206] = 8'h28;
s_mem_contents[14'h2207] = 8'ha9;
s_mem_contents[14'h2208] = 8'h00;
s_mem_contents[14'h2209] = 8'h48;
s_mem_contents[14'h220a] = 8'ha9;
s_mem_contents[14'h220b] = 8'h7f;
s_mem_contents[14'h220c] = 8'h28;
s_mem_contents[14'h220d] = 8'hd1;
s_mem_contents[14'h220e] = 8'h1a;
s_mem_contents[14'h220f] = 8'h08;
s_mem_contents[14'h2210] = 8'hc9;
s_mem_contents[14'h2211] = 8'h7f;
s_mem_contents[14'h2212] = 8'hd0;
s_mem_contents[14'h2213] = 8'hfe;
s_mem_contents[14'h2214] = 8'h68;
s_mem_contents[14'h2215] = 8'h48;
s_mem_contents[14'h2216] = 8'hc9;
s_mem_contents[14'h2217] = 8'h33;
s_mem_contents[14'h2218] = 8'hd0;
s_mem_contents[14'h2219] = 8'hfe;
s_mem_contents[14'h221a] = 8'h28;
s_mem_contents[14'h221b] = 8'ha9;
s_mem_contents[14'h221c] = 8'h00;
s_mem_contents[14'h221d] = 8'h48;
s_mem_contents[14'h221e] = 8'ha9;
s_mem_contents[14'h221f] = 8'h7e;
s_mem_contents[14'h2220] = 8'h28;
s_mem_contents[14'h2221] = 8'hd1;
s_mem_contents[14'h2222] = 8'h1a;
s_mem_contents[14'h2223] = 8'h08;
s_mem_contents[14'h2224] = 8'hc9;
s_mem_contents[14'h2225] = 8'h7e;
s_mem_contents[14'h2226] = 8'hd0;
s_mem_contents[14'h2227] = 8'hfe;
s_mem_contents[14'h2228] = 8'h68;
s_mem_contents[14'h2229] = 8'h48;
s_mem_contents[14'h222a] = 8'hc9;
s_mem_contents[14'h222b] = 8'hb0;
s_mem_contents[14'h222c] = 8'hd0;
s_mem_contents[14'h222d] = 8'hfe;
s_mem_contents[14'h222e] = 8'h28;
s_mem_contents[14'h222f] = 8'ha9;
s_mem_contents[14'h2230] = 8'hff;
s_mem_contents[14'h2231] = 8'h48;
s_mem_contents[14'h2232] = 8'ha9;
s_mem_contents[14'h2233] = 8'h80;
s_mem_contents[14'h2234] = 8'h28;
s_mem_contents[14'h2235] = 8'hd1;
s_mem_contents[14'h2236] = 8'h1a;
s_mem_contents[14'h2237] = 8'h08;
s_mem_contents[14'h2238] = 8'hc9;
s_mem_contents[14'h2239] = 8'h80;
s_mem_contents[14'h223a] = 8'hd0;
s_mem_contents[14'h223b] = 8'hfe;
s_mem_contents[14'h223c] = 8'h68;
s_mem_contents[14'h223d] = 8'h48;
s_mem_contents[14'h223e] = 8'hc9;
s_mem_contents[14'h223f] = 8'h7d;
s_mem_contents[14'h2240] = 8'hd0;
s_mem_contents[14'h2241] = 8'hfe;
s_mem_contents[14'h2242] = 8'h28;
s_mem_contents[14'h2243] = 8'ha9;
s_mem_contents[14'h2244] = 8'hff;
s_mem_contents[14'h2245] = 8'h48;
s_mem_contents[14'h2246] = 8'ha9;
s_mem_contents[14'h2247] = 8'h7f;
s_mem_contents[14'h2248] = 8'h28;
s_mem_contents[14'h2249] = 8'hd1;
s_mem_contents[14'h224a] = 8'h1a;
s_mem_contents[14'h224b] = 8'h08;
s_mem_contents[14'h224c] = 8'hc9;
s_mem_contents[14'h224d] = 8'h7f;
s_mem_contents[14'h224e] = 8'hd0;
s_mem_contents[14'h224f] = 8'hfe;
s_mem_contents[14'h2250] = 8'h68;
s_mem_contents[14'h2251] = 8'h48;
s_mem_contents[14'h2252] = 8'hc9;
s_mem_contents[14'h2253] = 8'h7f;
s_mem_contents[14'h2254] = 8'hd0;
s_mem_contents[14'h2255] = 8'hfe;
s_mem_contents[14'h2256] = 8'h28;
s_mem_contents[14'h2257] = 8'ha9;
s_mem_contents[14'h2258] = 8'hff;
s_mem_contents[14'h2259] = 8'h48;
s_mem_contents[14'h225a] = 8'ha9;
s_mem_contents[14'h225b] = 8'h7e;
s_mem_contents[14'h225c] = 8'h28;
s_mem_contents[14'h225d] = 8'hd1;
s_mem_contents[14'h225e] = 8'h1a;
s_mem_contents[14'h225f] = 8'h08;
s_mem_contents[14'h2260] = 8'hc9;
s_mem_contents[14'h2261] = 8'h7e;
s_mem_contents[14'h2262] = 8'hd0;
s_mem_contents[14'h2263] = 8'hfe;
s_mem_contents[14'h2264] = 8'h68;
s_mem_contents[14'h2265] = 8'h48;
s_mem_contents[14'h2266] = 8'hc9;
s_mem_contents[14'h2267] = 8'hfc;
s_mem_contents[14'h2268] = 8'hd0;
s_mem_contents[14'h2269] = 8'hfe;
s_mem_contents[14'h226a] = 8'h28;
s_mem_contents[14'h226b] = 8'had;
s_mem_contents[14'h226c] = 8'h00;
s_mem_contents[14'h226d] = 8'h02;
s_mem_contents[14'h226e] = 8'hc9;
s_mem_contents[14'h226f] = 8'h1c;
s_mem_contents[14'h2270] = 8'hd0;
s_mem_contents[14'h2271] = 8'hfe;
s_mem_contents[14'h2272] = 8'ha9;
s_mem_contents[14'h2273] = 8'h1d;
s_mem_contents[14'h2274] = 8'h8d;
s_mem_contents[14'h2275] = 8'h00;
s_mem_contents[14'h2276] = 8'h02;
s_mem_contents[14'h2277] = 8'ha2;
s_mem_contents[14'h2278] = 8'h03;
s_mem_contents[14'h2279] = 8'ha9;
s_mem_contents[14'h227a] = 8'h00;
s_mem_contents[14'h227b] = 8'h48;
s_mem_contents[14'h227c] = 8'hb5;
s_mem_contents[14'h227d] = 8'h09;
s_mem_contents[14'h227e] = 8'h28;
s_mem_contents[14'h227f] = 8'h0a;
s_mem_contents[14'h2280] = 8'h08;
s_mem_contents[14'h2281] = 8'hdd;
s_mem_contents[14'h2282] = 8'h20;
s_mem_contents[14'h2283] = 8'h02;
s_mem_contents[14'h2284] = 8'hd0;
s_mem_contents[14'h2285] = 8'hfe;
s_mem_contents[14'h2286] = 8'h68;
s_mem_contents[14'h2287] = 8'h49;
s_mem_contents[14'h2288] = 8'h30;
s_mem_contents[14'h2289] = 8'hdd;
s_mem_contents[14'h228a] = 8'h30;
s_mem_contents[14'h228b] = 8'h02;
s_mem_contents[14'h228c] = 8'hd0;
s_mem_contents[14'h228d] = 8'hfe;
s_mem_contents[14'h228e] = 8'hca;
s_mem_contents[14'h228f] = 8'h10;
s_mem_contents[14'h2290] = 8'he8;
s_mem_contents[14'h2291] = 8'ha2;
s_mem_contents[14'h2292] = 8'h03;
s_mem_contents[14'h2293] = 8'ha9;
s_mem_contents[14'h2294] = 8'hff;
s_mem_contents[14'h2295] = 8'h48;
s_mem_contents[14'h2296] = 8'hb5;
s_mem_contents[14'h2297] = 8'h09;
s_mem_contents[14'h2298] = 8'h28;
s_mem_contents[14'h2299] = 8'h0a;
s_mem_contents[14'h229a] = 8'h08;
s_mem_contents[14'h229b] = 8'hdd;
s_mem_contents[14'h229c] = 8'h20;
s_mem_contents[14'h229d] = 8'h02;
s_mem_contents[14'h229e] = 8'hd0;
s_mem_contents[14'h229f] = 8'hfe;
s_mem_contents[14'h22a0] = 8'h68;
s_mem_contents[14'h22a1] = 8'h49;
s_mem_contents[14'h22a2] = 8'h7c;
s_mem_contents[14'h22a3] = 8'hdd;
s_mem_contents[14'h22a4] = 8'h30;
s_mem_contents[14'h22a5] = 8'h02;
s_mem_contents[14'h22a6] = 8'hd0;
s_mem_contents[14'h22a7] = 8'hfe;
s_mem_contents[14'h22a8] = 8'hca;
s_mem_contents[14'h22a9] = 8'h10;
s_mem_contents[14'h22aa] = 8'he8;
s_mem_contents[14'h22ab] = 8'ha2;
s_mem_contents[14'h22ac] = 8'h03;
s_mem_contents[14'h22ad] = 8'ha9;
s_mem_contents[14'h22ae] = 8'h00;
s_mem_contents[14'h22af] = 8'h48;
s_mem_contents[14'h22b0] = 8'hb5;
s_mem_contents[14'h22b1] = 8'h09;
s_mem_contents[14'h22b2] = 8'h28;
s_mem_contents[14'h22b3] = 8'h4a;
s_mem_contents[14'h22b4] = 8'h08;
s_mem_contents[14'h22b5] = 8'hdd;
s_mem_contents[14'h22b6] = 8'h28;
s_mem_contents[14'h22b7] = 8'h02;
s_mem_contents[14'h22b8] = 8'hd0;
s_mem_contents[14'h22b9] = 8'hfe;
s_mem_contents[14'h22ba] = 8'h68;
s_mem_contents[14'h22bb] = 8'h49;
s_mem_contents[14'h22bc] = 8'h30;
s_mem_contents[14'h22bd] = 8'hdd;
s_mem_contents[14'h22be] = 8'h38;
s_mem_contents[14'h22bf] = 8'h02;
s_mem_contents[14'h22c0] = 8'hd0;
s_mem_contents[14'h22c1] = 8'hfe;
s_mem_contents[14'h22c2] = 8'hca;
s_mem_contents[14'h22c3] = 8'h10;
s_mem_contents[14'h22c4] = 8'he8;
s_mem_contents[14'h22c5] = 8'ha2;
s_mem_contents[14'h22c6] = 8'h03;
s_mem_contents[14'h22c7] = 8'ha9;
s_mem_contents[14'h22c8] = 8'hff;
s_mem_contents[14'h22c9] = 8'h48;
s_mem_contents[14'h22ca] = 8'hb5;
s_mem_contents[14'h22cb] = 8'h09;
s_mem_contents[14'h22cc] = 8'h28;
s_mem_contents[14'h22cd] = 8'h4a;
s_mem_contents[14'h22ce] = 8'h08;
s_mem_contents[14'h22cf] = 8'hdd;
s_mem_contents[14'h22d0] = 8'h28;
s_mem_contents[14'h22d1] = 8'h02;
s_mem_contents[14'h22d2] = 8'hd0;
s_mem_contents[14'h22d3] = 8'hfe;
s_mem_contents[14'h22d4] = 8'h68;
s_mem_contents[14'h22d5] = 8'h49;
s_mem_contents[14'h22d6] = 8'h7c;
s_mem_contents[14'h22d7] = 8'hdd;
s_mem_contents[14'h22d8] = 8'h38;
s_mem_contents[14'h22d9] = 8'h02;
s_mem_contents[14'h22da] = 8'hd0;
s_mem_contents[14'h22db] = 8'hfe;
s_mem_contents[14'h22dc] = 8'hca;
s_mem_contents[14'h22dd] = 8'h10;
s_mem_contents[14'h22de] = 8'he8;
s_mem_contents[14'h22df] = 8'ha2;
s_mem_contents[14'h22e0] = 8'h03;
s_mem_contents[14'h22e1] = 8'ha9;
s_mem_contents[14'h22e2] = 8'h00;
s_mem_contents[14'h22e3] = 8'h48;
s_mem_contents[14'h22e4] = 8'hb5;
s_mem_contents[14'h22e5] = 8'h09;
s_mem_contents[14'h22e6] = 8'h28;
s_mem_contents[14'h22e7] = 8'h2a;
s_mem_contents[14'h22e8] = 8'h08;
s_mem_contents[14'h22e9] = 8'hdd;
s_mem_contents[14'h22ea] = 8'h20;
s_mem_contents[14'h22eb] = 8'h02;
s_mem_contents[14'h22ec] = 8'hd0;
s_mem_contents[14'h22ed] = 8'hfe;
s_mem_contents[14'h22ee] = 8'h68;
s_mem_contents[14'h22ef] = 8'h49;
s_mem_contents[14'h22f0] = 8'h30;
s_mem_contents[14'h22f1] = 8'hdd;
s_mem_contents[14'h22f2] = 8'h30;
s_mem_contents[14'h22f3] = 8'h02;
s_mem_contents[14'h22f4] = 8'hd0;
s_mem_contents[14'h22f5] = 8'hfe;
s_mem_contents[14'h22f6] = 8'hca;
s_mem_contents[14'h22f7] = 8'h10;
s_mem_contents[14'h22f8] = 8'he8;
s_mem_contents[14'h22f9] = 8'ha2;
s_mem_contents[14'h22fa] = 8'h03;
s_mem_contents[14'h22fb] = 8'ha9;
s_mem_contents[14'h22fc] = 8'hfe;
s_mem_contents[14'h22fd] = 8'h48;
s_mem_contents[14'h22fe] = 8'hb5;
s_mem_contents[14'h22ff] = 8'h09;
s_mem_contents[14'h2300] = 8'h28;
s_mem_contents[14'h2301] = 8'h2a;
s_mem_contents[14'h2302] = 8'h08;
s_mem_contents[14'h2303] = 8'hdd;
s_mem_contents[14'h2304] = 8'h20;
s_mem_contents[14'h2305] = 8'h02;
s_mem_contents[14'h2306] = 8'hd0;
s_mem_contents[14'h2307] = 8'hfe;
s_mem_contents[14'h2308] = 8'h68;
s_mem_contents[14'h2309] = 8'h49;
s_mem_contents[14'h230a] = 8'h7c;
s_mem_contents[14'h230b] = 8'hdd;
s_mem_contents[14'h230c] = 8'h30;
s_mem_contents[14'h230d] = 8'h02;
s_mem_contents[14'h230e] = 8'hd0;
s_mem_contents[14'h230f] = 8'hfe;
s_mem_contents[14'h2310] = 8'hca;
s_mem_contents[14'h2311] = 8'h10;
s_mem_contents[14'h2312] = 8'he8;
s_mem_contents[14'h2313] = 8'ha2;
s_mem_contents[14'h2314] = 8'h03;
s_mem_contents[14'h2315] = 8'ha9;
s_mem_contents[14'h2316] = 8'h01;
s_mem_contents[14'h2317] = 8'h48;
s_mem_contents[14'h2318] = 8'hb5;
s_mem_contents[14'h2319] = 8'h09;
s_mem_contents[14'h231a] = 8'h28;
s_mem_contents[14'h231b] = 8'h2a;
s_mem_contents[14'h231c] = 8'h08;
s_mem_contents[14'h231d] = 8'hdd;
s_mem_contents[14'h231e] = 8'h24;
s_mem_contents[14'h231f] = 8'h02;
s_mem_contents[14'h2320] = 8'hd0;
s_mem_contents[14'h2321] = 8'hfe;
s_mem_contents[14'h2322] = 8'h68;
s_mem_contents[14'h2323] = 8'h49;
s_mem_contents[14'h2324] = 8'h30;
s_mem_contents[14'h2325] = 8'hdd;
s_mem_contents[14'h2326] = 8'h34;
s_mem_contents[14'h2327] = 8'h02;
s_mem_contents[14'h2328] = 8'hd0;
s_mem_contents[14'h2329] = 8'hfe;
s_mem_contents[14'h232a] = 8'hca;
s_mem_contents[14'h232b] = 8'h10;
s_mem_contents[14'h232c] = 8'he8;
s_mem_contents[14'h232d] = 8'ha2;
s_mem_contents[14'h232e] = 8'h03;
s_mem_contents[14'h232f] = 8'ha9;
s_mem_contents[14'h2330] = 8'hff;
s_mem_contents[14'h2331] = 8'h48;
s_mem_contents[14'h2332] = 8'hb5;
s_mem_contents[14'h2333] = 8'h09;
s_mem_contents[14'h2334] = 8'h28;
s_mem_contents[14'h2335] = 8'h2a;
s_mem_contents[14'h2336] = 8'h08;
s_mem_contents[14'h2337] = 8'hdd;
s_mem_contents[14'h2338] = 8'h24;
s_mem_contents[14'h2339] = 8'h02;
s_mem_contents[14'h233a] = 8'hd0;
s_mem_contents[14'h233b] = 8'hfe;
s_mem_contents[14'h233c] = 8'h68;
s_mem_contents[14'h233d] = 8'h49;
s_mem_contents[14'h233e] = 8'h7c;
s_mem_contents[14'h233f] = 8'hdd;
s_mem_contents[14'h2340] = 8'h34;
s_mem_contents[14'h2341] = 8'h02;
s_mem_contents[14'h2342] = 8'hd0;
s_mem_contents[14'h2343] = 8'hfe;
s_mem_contents[14'h2344] = 8'hca;
s_mem_contents[14'h2345] = 8'h10;
s_mem_contents[14'h2346] = 8'he8;
s_mem_contents[14'h2347] = 8'ha2;
s_mem_contents[14'h2348] = 8'h03;
s_mem_contents[14'h2349] = 8'ha9;
s_mem_contents[14'h234a] = 8'h00;
s_mem_contents[14'h234b] = 8'h48;
s_mem_contents[14'h234c] = 8'hb5;
s_mem_contents[14'h234d] = 8'h09;
s_mem_contents[14'h234e] = 8'h28;
s_mem_contents[14'h234f] = 8'h6a;
s_mem_contents[14'h2350] = 8'h08;
s_mem_contents[14'h2351] = 8'hdd;
s_mem_contents[14'h2352] = 8'h28;
s_mem_contents[14'h2353] = 8'h02;
s_mem_contents[14'h2354] = 8'hd0;
s_mem_contents[14'h2355] = 8'hfe;
s_mem_contents[14'h2356] = 8'h68;
s_mem_contents[14'h2357] = 8'h49;
s_mem_contents[14'h2358] = 8'h30;
s_mem_contents[14'h2359] = 8'hdd;
s_mem_contents[14'h235a] = 8'h38;
s_mem_contents[14'h235b] = 8'h02;
s_mem_contents[14'h235c] = 8'hd0;
s_mem_contents[14'h235d] = 8'hfe;
s_mem_contents[14'h235e] = 8'hca;
s_mem_contents[14'h235f] = 8'h10;
s_mem_contents[14'h2360] = 8'he8;
s_mem_contents[14'h2361] = 8'ha2;
s_mem_contents[14'h2362] = 8'h03;
s_mem_contents[14'h2363] = 8'ha9;
s_mem_contents[14'h2364] = 8'hfe;
s_mem_contents[14'h2365] = 8'h48;
s_mem_contents[14'h2366] = 8'hb5;
s_mem_contents[14'h2367] = 8'h09;
s_mem_contents[14'h2368] = 8'h28;
s_mem_contents[14'h2369] = 8'h6a;
s_mem_contents[14'h236a] = 8'h08;
s_mem_contents[14'h236b] = 8'hdd;
s_mem_contents[14'h236c] = 8'h28;
s_mem_contents[14'h236d] = 8'h02;
s_mem_contents[14'h236e] = 8'hd0;
s_mem_contents[14'h236f] = 8'hfe;
s_mem_contents[14'h2370] = 8'h68;
s_mem_contents[14'h2371] = 8'h49;
s_mem_contents[14'h2372] = 8'h7c;
s_mem_contents[14'h2373] = 8'hdd;
s_mem_contents[14'h2374] = 8'h38;
s_mem_contents[14'h2375] = 8'h02;
s_mem_contents[14'h2376] = 8'hd0;
s_mem_contents[14'h2377] = 8'hfe;
s_mem_contents[14'h2378] = 8'hca;
s_mem_contents[14'h2379] = 8'h10;
s_mem_contents[14'h237a] = 8'he8;
s_mem_contents[14'h237b] = 8'ha2;
s_mem_contents[14'h237c] = 8'h03;
s_mem_contents[14'h237d] = 8'ha9;
s_mem_contents[14'h237e] = 8'h01;
s_mem_contents[14'h237f] = 8'h48;
s_mem_contents[14'h2380] = 8'hb5;
s_mem_contents[14'h2381] = 8'h09;
s_mem_contents[14'h2382] = 8'h28;
s_mem_contents[14'h2383] = 8'h6a;
s_mem_contents[14'h2384] = 8'h08;
s_mem_contents[14'h2385] = 8'hdd;
s_mem_contents[14'h2386] = 8'h2c;
s_mem_contents[14'h2387] = 8'h02;
s_mem_contents[14'h2388] = 8'hd0;
s_mem_contents[14'h2389] = 8'hfe;
s_mem_contents[14'h238a] = 8'h68;
s_mem_contents[14'h238b] = 8'h49;
s_mem_contents[14'h238c] = 8'h30;
s_mem_contents[14'h238d] = 8'hdd;
s_mem_contents[14'h238e] = 8'h3c;
s_mem_contents[14'h238f] = 8'h02;
s_mem_contents[14'h2390] = 8'hd0;
s_mem_contents[14'h2391] = 8'hfe;
s_mem_contents[14'h2392] = 8'hca;
s_mem_contents[14'h2393] = 8'h10;
s_mem_contents[14'h2394] = 8'he8;
s_mem_contents[14'h2395] = 8'ha2;
s_mem_contents[14'h2396] = 8'h03;
s_mem_contents[14'h2397] = 8'ha9;
s_mem_contents[14'h2398] = 8'hff;
s_mem_contents[14'h2399] = 8'h48;
s_mem_contents[14'h239a] = 8'hb5;
s_mem_contents[14'h239b] = 8'h09;
s_mem_contents[14'h239c] = 8'h28;
s_mem_contents[14'h239d] = 8'h6a;
s_mem_contents[14'h239e] = 8'h08;
s_mem_contents[14'h239f] = 8'hdd;
s_mem_contents[14'h23a0] = 8'h2c;
s_mem_contents[14'h23a1] = 8'h02;
s_mem_contents[14'h23a2] = 8'hd0;
s_mem_contents[14'h23a3] = 8'hfe;
s_mem_contents[14'h23a4] = 8'h68;
s_mem_contents[14'h23a5] = 8'h49;
s_mem_contents[14'h23a6] = 8'h7c;
s_mem_contents[14'h23a7] = 8'hdd;
s_mem_contents[14'h23a8] = 8'h3c;
s_mem_contents[14'h23a9] = 8'h02;
s_mem_contents[14'h23aa] = 8'hd0;
s_mem_contents[14'h23ab] = 8'hfe;
s_mem_contents[14'h23ac] = 8'hca;
s_mem_contents[14'h23ad] = 8'h10;
s_mem_contents[14'h23ae] = 8'he8;
s_mem_contents[14'h23af] = 8'had;
s_mem_contents[14'h23b0] = 8'h00;
s_mem_contents[14'h23b1] = 8'h02;
s_mem_contents[14'h23b2] = 8'hc9;
s_mem_contents[14'h23b3] = 8'h1d;
s_mem_contents[14'h23b4] = 8'hd0;
s_mem_contents[14'h23b5] = 8'hfe;
s_mem_contents[14'h23b6] = 8'ha9;
s_mem_contents[14'h23b7] = 8'h1e;
s_mem_contents[14'h23b8] = 8'h8d;
s_mem_contents[14'h23b9] = 8'h00;
s_mem_contents[14'h23ba] = 8'h02;
s_mem_contents[14'h23bb] = 8'ha2;
s_mem_contents[14'h23bc] = 8'h03;
s_mem_contents[14'h23bd] = 8'ha9;
s_mem_contents[14'h23be] = 8'h00;
s_mem_contents[14'h23bf] = 8'h48;
s_mem_contents[14'h23c0] = 8'hb5;
s_mem_contents[14'h23c1] = 8'h09;
s_mem_contents[14'h23c2] = 8'h85;
s_mem_contents[14'h23c3] = 8'h02;
s_mem_contents[14'h23c4] = 8'h28;
s_mem_contents[14'h23c5] = 8'h06;
s_mem_contents[14'h23c6] = 8'h02;
s_mem_contents[14'h23c7] = 8'h08;
s_mem_contents[14'h23c8] = 8'ha5;
s_mem_contents[14'h23c9] = 8'h02;
s_mem_contents[14'h23ca] = 8'hdd;
s_mem_contents[14'h23cb] = 8'h20;
s_mem_contents[14'h23cc] = 8'h02;
s_mem_contents[14'h23cd] = 8'hd0;
s_mem_contents[14'h23ce] = 8'hfe;
s_mem_contents[14'h23cf] = 8'h68;
s_mem_contents[14'h23d0] = 8'h49;
s_mem_contents[14'h23d1] = 8'h30;
s_mem_contents[14'h23d2] = 8'hdd;
s_mem_contents[14'h23d3] = 8'h30;
s_mem_contents[14'h23d4] = 8'h02;
s_mem_contents[14'h23d5] = 8'hd0;
s_mem_contents[14'h23d6] = 8'hfe;
s_mem_contents[14'h23d7] = 8'hca;
s_mem_contents[14'h23d8] = 8'h10;
s_mem_contents[14'h23d9] = 8'he3;
s_mem_contents[14'h23da] = 8'ha2;
s_mem_contents[14'h23db] = 8'h03;
s_mem_contents[14'h23dc] = 8'ha9;
s_mem_contents[14'h23dd] = 8'hff;
s_mem_contents[14'h23de] = 8'h48;
s_mem_contents[14'h23df] = 8'hb5;
s_mem_contents[14'h23e0] = 8'h09;
s_mem_contents[14'h23e1] = 8'h85;
s_mem_contents[14'h23e2] = 8'h02;
s_mem_contents[14'h23e3] = 8'h28;
s_mem_contents[14'h23e4] = 8'h06;
s_mem_contents[14'h23e5] = 8'h02;
s_mem_contents[14'h23e6] = 8'h08;
s_mem_contents[14'h23e7] = 8'ha5;
s_mem_contents[14'h23e8] = 8'h02;
s_mem_contents[14'h23e9] = 8'hdd;
s_mem_contents[14'h23ea] = 8'h20;
s_mem_contents[14'h23eb] = 8'h02;
s_mem_contents[14'h23ec] = 8'hd0;
s_mem_contents[14'h23ed] = 8'hfe;
s_mem_contents[14'h23ee] = 8'h68;
s_mem_contents[14'h23ef] = 8'h49;
s_mem_contents[14'h23f0] = 8'h7c;
s_mem_contents[14'h23f1] = 8'hdd;
s_mem_contents[14'h23f2] = 8'h30;
s_mem_contents[14'h23f3] = 8'h02;
s_mem_contents[14'h23f4] = 8'hd0;
s_mem_contents[14'h23f5] = 8'hfe;
s_mem_contents[14'h23f6] = 8'hca;
s_mem_contents[14'h23f7] = 8'h10;
s_mem_contents[14'h23f8] = 8'he3;
s_mem_contents[14'h23f9] = 8'ha2;
s_mem_contents[14'h23fa] = 8'h03;
s_mem_contents[14'h23fb] = 8'ha9;
s_mem_contents[14'h23fc] = 8'h00;
s_mem_contents[14'h23fd] = 8'h48;
s_mem_contents[14'h23fe] = 8'hb5;
s_mem_contents[14'h23ff] = 8'h09;
s_mem_contents[14'h2400] = 8'h85;
s_mem_contents[14'h2401] = 8'h02;
s_mem_contents[14'h2402] = 8'h28;
s_mem_contents[14'h2403] = 8'h46;
s_mem_contents[14'h2404] = 8'h02;
s_mem_contents[14'h2405] = 8'h08;
s_mem_contents[14'h2406] = 8'ha5;
s_mem_contents[14'h2407] = 8'h02;
s_mem_contents[14'h2408] = 8'hdd;
s_mem_contents[14'h2409] = 8'h28;
s_mem_contents[14'h240a] = 8'h02;
s_mem_contents[14'h240b] = 8'hd0;
s_mem_contents[14'h240c] = 8'hfe;
s_mem_contents[14'h240d] = 8'h68;
s_mem_contents[14'h240e] = 8'h49;
s_mem_contents[14'h240f] = 8'h30;
s_mem_contents[14'h2410] = 8'hdd;
s_mem_contents[14'h2411] = 8'h38;
s_mem_contents[14'h2412] = 8'h02;
s_mem_contents[14'h2413] = 8'hd0;
s_mem_contents[14'h2414] = 8'hfe;
s_mem_contents[14'h2415] = 8'hca;
s_mem_contents[14'h2416] = 8'h10;
s_mem_contents[14'h2417] = 8'he3;
s_mem_contents[14'h2418] = 8'ha2;
s_mem_contents[14'h2419] = 8'h03;
s_mem_contents[14'h241a] = 8'ha9;
s_mem_contents[14'h241b] = 8'hff;
s_mem_contents[14'h241c] = 8'h48;
s_mem_contents[14'h241d] = 8'hb5;
s_mem_contents[14'h241e] = 8'h09;
s_mem_contents[14'h241f] = 8'h85;
s_mem_contents[14'h2420] = 8'h02;
s_mem_contents[14'h2421] = 8'h28;
s_mem_contents[14'h2422] = 8'h46;
s_mem_contents[14'h2423] = 8'h02;
s_mem_contents[14'h2424] = 8'h08;
s_mem_contents[14'h2425] = 8'ha5;
s_mem_contents[14'h2426] = 8'h02;
s_mem_contents[14'h2427] = 8'hdd;
s_mem_contents[14'h2428] = 8'h28;
s_mem_contents[14'h2429] = 8'h02;
s_mem_contents[14'h242a] = 8'hd0;
s_mem_contents[14'h242b] = 8'hfe;
s_mem_contents[14'h242c] = 8'h68;
s_mem_contents[14'h242d] = 8'h49;
s_mem_contents[14'h242e] = 8'h7c;
s_mem_contents[14'h242f] = 8'hdd;
s_mem_contents[14'h2430] = 8'h38;
s_mem_contents[14'h2431] = 8'h02;
s_mem_contents[14'h2432] = 8'hd0;
s_mem_contents[14'h2433] = 8'hfe;
s_mem_contents[14'h2434] = 8'hca;
s_mem_contents[14'h2435] = 8'h10;
s_mem_contents[14'h2436] = 8'he3;
s_mem_contents[14'h2437] = 8'ha2;
s_mem_contents[14'h2438] = 8'h03;
s_mem_contents[14'h2439] = 8'ha9;
s_mem_contents[14'h243a] = 8'h00;
s_mem_contents[14'h243b] = 8'h48;
s_mem_contents[14'h243c] = 8'hb5;
s_mem_contents[14'h243d] = 8'h09;
s_mem_contents[14'h243e] = 8'h85;
s_mem_contents[14'h243f] = 8'h02;
s_mem_contents[14'h2440] = 8'h28;
s_mem_contents[14'h2441] = 8'h26;
s_mem_contents[14'h2442] = 8'h02;
s_mem_contents[14'h2443] = 8'h08;
s_mem_contents[14'h2444] = 8'ha5;
s_mem_contents[14'h2445] = 8'h02;
s_mem_contents[14'h2446] = 8'hdd;
s_mem_contents[14'h2447] = 8'h20;
s_mem_contents[14'h2448] = 8'h02;
s_mem_contents[14'h2449] = 8'hd0;
s_mem_contents[14'h244a] = 8'hfe;
s_mem_contents[14'h244b] = 8'h68;
s_mem_contents[14'h244c] = 8'h49;
s_mem_contents[14'h244d] = 8'h30;
s_mem_contents[14'h244e] = 8'hdd;
s_mem_contents[14'h244f] = 8'h30;
s_mem_contents[14'h2450] = 8'h02;
s_mem_contents[14'h2451] = 8'hd0;
s_mem_contents[14'h2452] = 8'hfe;
s_mem_contents[14'h2453] = 8'hca;
s_mem_contents[14'h2454] = 8'h10;
s_mem_contents[14'h2455] = 8'he3;
s_mem_contents[14'h2456] = 8'ha2;
s_mem_contents[14'h2457] = 8'h03;
s_mem_contents[14'h2458] = 8'ha9;
s_mem_contents[14'h2459] = 8'hfe;
s_mem_contents[14'h245a] = 8'h48;
s_mem_contents[14'h245b] = 8'hb5;
s_mem_contents[14'h245c] = 8'h09;
s_mem_contents[14'h245d] = 8'h85;
s_mem_contents[14'h245e] = 8'h02;
s_mem_contents[14'h245f] = 8'h28;
s_mem_contents[14'h2460] = 8'h26;
s_mem_contents[14'h2461] = 8'h02;
s_mem_contents[14'h2462] = 8'h08;
s_mem_contents[14'h2463] = 8'ha5;
s_mem_contents[14'h2464] = 8'h02;
s_mem_contents[14'h2465] = 8'hdd;
s_mem_contents[14'h2466] = 8'h20;
s_mem_contents[14'h2467] = 8'h02;
s_mem_contents[14'h2468] = 8'hd0;
s_mem_contents[14'h2469] = 8'hfe;
s_mem_contents[14'h246a] = 8'h68;
s_mem_contents[14'h246b] = 8'h49;
s_mem_contents[14'h246c] = 8'h7c;
s_mem_contents[14'h246d] = 8'hdd;
s_mem_contents[14'h246e] = 8'h30;
s_mem_contents[14'h246f] = 8'h02;
s_mem_contents[14'h2470] = 8'hd0;
s_mem_contents[14'h2471] = 8'hfe;
s_mem_contents[14'h2472] = 8'hca;
s_mem_contents[14'h2473] = 8'h10;
s_mem_contents[14'h2474] = 8'he3;
s_mem_contents[14'h2475] = 8'ha2;
s_mem_contents[14'h2476] = 8'h03;
s_mem_contents[14'h2477] = 8'ha9;
s_mem_contents[14'h2478] = 8'h01;
s_mem_contents[14'h2479] = 8'h48;
s_mem_contents[14'h247a] = 8'hb5;
s_mem_contents[14'h247b] = 8'h09;
s_mem_contents[14'h247c] = 8'h85;
s_mem_contents[14'h247d] = 8'h02;
s_mem_contents[14'h247e] = 8'h28;
s_mem_contents[14'h247f] = 8'h26;
s_mem_contents[14'h2480] = 8'h02;
s_mem_contents[14'h2481] = 8'h08;
s_mem_contents[14'h2482] = 8'ha5;
s_mem_contents[14'h2483] = 8'h02;
s_mem_contents[14'h2484] = 8'hdd;
s_mem_contents[14'h2485] = 8'h24;
s_mem_contents[14'h2486] = 8'h02;
s_mem_contents[14'h2487] = 8'hd0;
s_mem_contents[14'h2488] = 8'hfe;
s_mem_contents[14'h2489] = 8'h68;
s_mem_contents[14'h248a] = 8'h49;
s_mem_contents[14'h248b] = 8'h30;
s_mem_contents[14'h248c] = 8'hdd;
s_mem_contents[14'h248d] = 8'h34;
s_mem_contents[14'h248e] = 8'h02;
s_mem_contents[14'h248f] = 8'hd0;
s_mem_contents[14'h2490] = 8'hfe;
s_mem_contents[14'h2491] = 8'hca;
s_mem_contents[14'h2492] = 8'h10;
s_mem_contents[14'h2493] = 8'he3;
s_mem_contents[14'h2494] = 8'ha2;
s_mem_contents[14'h2495] = 8'h03;
s_mem_contents[14'h2496] = 8'ha9;
s_mem_contents[14'h2497] = 8'hff;
s_mem_contents[14'h2498] = 8'h48;
s_mem_contents[14'h2499] = 8'hb5;
s_mem_contents[14'h249a] = 8'h09;
s_mem_contents[14'h249b] = 8'h85;
s_mem_contents[14'h249c] = 8'h02;
s_mem_contents[14'h249d] = 8'h28;
s_mem_contents[14'h249e] = 8'h26;
s_mem_contents[14'h249f] = 8'h02;
s_mem_contents[14'h24a0] = 8'h08;
s_mem_contents[14'h24a1] = 8'ha5;
s_mem_contents[14'h24a2] = 8'h02;
s_mem_contents[14'h24a3] = 8'hdd;
s_mem_contents[14'h24a4] = 8'h24;
s_mem_contents[14'h24a5] = 8'h02;
s_mem_contents[14'h24a6] = 8'hd0;
s_mem_contents[14'h24a7] = 8'hfe;
s_mem_contents[14'h24a8] = 8'h68;
s_mem_contents[14'h24a9] = 8'h49;
s_mem_contents[14'h24aa] = 8'h7c;
s_mem_contents[14'h24ab] = 8'hdd;
s_mem_contents[14'h24ac] = 8'h34;
s_mem_contents[14'h24ad] = 8'h02;
s_mem_contents[14'h24ae] = 8'hd0;
s_mem_contents[14'h24af] = 8'hfe;
s_mem_contents[14'h24b0] = 8'hca;
s_mem_contents[14'h24b1] = 8'h10;
s_mem_contents[14'h24b2] = 8'he3;
s_mem_contents[14'h24b3] = 8'ha2;
s_mem_contents[14'h24b4] = 8'h03;
s_mem_contents[14'h24b5] = 8'ha9;
s_mem_contents[14'h24b6] = 8'h00;
s_mem_contents[14'h24b7] = 8'h48;
s_mem_contents[14'h24b8] = 8'hb5;
s_mem_contents[14'h24b9] = 8'h09;
s_mem_contents[14'h24ba] = 8'h85;
s_mem_contents[14'h24bb] = 8'h02;
s_mem_contents[14'h24bc] = 8'h28;
s_mem_contents[14'h24bd] = 8'h66;
s_mem_contents[14'h24be] = 8'h02;
s_mem_contents[14'h24bf] = 8'h08;
s_mem_contents[14'h24c0] = 8'ha5;
s_mem_contents[14'h24c1] = 8'h02;
s_mem_contents[14'h24c2] = 8'hdd;
s_mem_contents[14'h24c3] = 8'h28;
s_mem_contents[14'h24c4] = 8'h02;
s_mem_contents[14'h24c5] = 8'hd0;
s_mem_contents[14'h24c6] = 8'hfe;
s_mem_contents[14'h24c7] = 8'h68;
s_mem_contents[14'h24c8] = 8'h49;
s_mem_contents[14'h24c9] = 8'h30;
s_mem_contents[14'h24ca] = 8'hdd;
s_mem_contents[14'h24cb] = 8'h38;
s_mem_contents[14'h24cc] = 8'h02;
s_mem_contents[14'h24cd] = 8'hd0;
s_mem_contents[14'h24ce] = 8'hfe;
s_mem_contents[14'h24cf] = 8'hca;
s_mem_contents[14'h24d0] = 8'h10;
s_mem_contents[14'h24d1] = 8'he3;
s_mem_contents[14'h24d2] = 8'ha2;
s_mem_contents[14'h24d3] = 8'h03;
s_mem_contents[14'h24d4] = 8'ha9;
s_mem_contents[14'h24d5] = 8'hfe;
s_mem_contents[14'h24d6] = 8'h48;
s_mem_contents[14'h24d7] = 8'hb5;
s_mem_contents[14'h24d8] = 8'h09;
s_mem_contents[14'h24d9] = 8'h85;
s_mem_contents[14'h24da] = 8'h02;
s_mem_contents[14'h24db] = 8'h28;
s_mem_contents[14'h24dc] = 8'h66;
s_mem_contents[14'h24dd] = 8'h02;
s_mem_contents[14'h24de] = 8'h08;
s_mem_contents[14'h24df] = 8'ha5;
s_mem_contents[14'h24e0] = 8'h02;
s_mem_contents[14'h24e1] = 8'hdd;
s_mem_contents[14'h24e2] = 8'h28;
s_mem_contents[14'h24e3] = 8'h02;
s_mem_contents[14'h24e4] = 8'hd0;
s_mem_contents[14'h24e5] = 8'hfe;
s_mem_contents[14'h24e6] = 8'h68;
s_mem_contents[14'h24e7] = 8'h49;
s_mem_contents[14'h24e8] = 8'h7c;
s_mem_contents[14'h24e9] = 8'hdd;
s_mem_contents[14'h24ea] = 8'h38;
s_mem_contents[14'h24eb] = 8'h02;
s_mem_contents[14'h24ec] = 8'hd0;
s_mem_contents[14'h24ed] = 8'hfe;
s_mem_contents[14'h24ee] = 8'hca;
s_mem_contents[14'h24ef] = 8'h10;
s_mem_contents[14'h24f0] = 8'he3;
s_mem_contents[14'h24f1] = 8'ha2;
s_mem_contents[14'h24f2] = 8'h03;
s_mem_contents[14'h24f3] = 8'ha9;
s_mem_contents[14'h24f4] = 8'h01;
s_mem_contents[14'h24f5] = 8'h48;
s_mem_contents[14'h24f6] = 8'hb5;
s_mem_contents[14'h24f7] = 8'h09;
s_mem_contents[14'h24f8] = 8'h85;
s_mem_contents[14'h24f9] = 8'h02;
s_mem_contents[14'h24fa] = 8'h28;
s_mem_contents[14'h24fb] = 8'h66;
s_mem_contents[14'h24fc] = 8'h02;
s_mem_contents[14'h24fd] = 8'h08;
s_mem_contents[14'h24fe] = 8'ha5;
s_mem_contents[14'h24ff] = 8'h02;
s_mem_contents[14'h2500] = 8'hdd;
s_mem_contents[14'h2501] = 8'h2c;
s_mem_contents[14'h2502] = 8'h02;
s_mem_contents[14'h2503] = 8'hd0;
s_mem_contents[14'h2504] = 8'hfe;
s_mem_contents[14'h2505] = 8'h68;
s_mem_contents[14'h2506] = 8'h49;
s_mem_contents[14'h2507] = 8'h30;
s_mem_contents[14'h2508] = 8'hdd;
s_mem_contents[14'h2509] = 8'h3c;
s_mem_contents[14'h250a] = 8'h02;
s_mem_contents[14'h250b] = 8'hd0;
s_mem_contents[14'h250c] = 8'hfe;
s_mem_contents[14'h250d] = 8'hca;
s_mem_contents[14'h250e] = 8'h10;
s_mem_contents[14'h250f] = 8'he3;
s_mem_contents[14'h2510] = 8'ha2;
s_mem_contents[14'h2511] = 8'h03;
s_mem_contents[14'h2512] = 8'ha9;
s_mem_contents[14'h2513] = 8'hff;
s_mem_contents[14'h2514] = 8'h48;
s_mem_contents[14'h2515] = 8'hb5;
s_mem_contents[14'h2516] = 8'h09;
s_mem_contents[14'h2517] = 8'h85;
s_mem_contents[14'h2518] = 8'h02;
s_mem_contents[14'h2519] = 8'h28;
s_mem_contents[14'h251a] = 8'h66;
s_mem_contents[14'h251b] = 8'h02;
s_mem_contents[14'h251c] = 8'h08;
s_mem_contents[14'h251d] = 8'ha5;
s_mem_contents[14'h251e] = 8'h02;
s_mem_contents[14'h251f] = 8'hdd;
s_mem_contents[14'h2520] = 8'h2c;
s_mem_contents[14'h2521] = 8'h02;
s_mem_contents[14'h2522] = 8'hd0;
s_mem_contents[14'h2523] = 8'hfe;
s_mem_contents[14'h2524] = 8'h68;
s_mem_contents[14'h2525] = 8'h49;
s_mem_contents[14'h2526] = 8'h7c;
s_mem_contents[14'h2527] = 8'hdd;
s_mem_contents[14'h2528] = 8'h3c;
s_mem_contents[14'h2529] = 8'h02;
s_mem_contents[14'h252a] = 8'hd0;
s_mem_contents[14'h252b] = 8'hfe;
s_mem_contents[14'h252c] = 8'hca;
s_mem_contents[14'h252d] = 8'h10;
s_mem_contents[14'h252e] = 8'he3;
s_mem_contents[14'h252f] = 8'had;
s_mem_contents[14'h2530] = 8'h00;
s_mem_contents[14'h2531] = 8'h02;
s_mem_contents[14'h2532] = 8'hc9;
s_mem_contents[14'h2533] = 8'h1e;
s_mem_contents[14'h2534] = 8'hd0;
s_mem_contents[14'h2535] = 8'hfe;
s_mem_contents[14'h2536] = 8'ha9;
s_mem_contents[14'h2537] = 8'h1f;
s_mem_contents[14'h2538] = 8'h8d;
s_mem_contents[14'h2539] = 8'h00;
s_mem_contents[14'h253a] = 8'h02;
s_mem_contents[14'h253b] = 8'ha2;
s_mem_contents[14'h253c] = 8'h03;
s_mem_contents[14'h253d] = 8'ha9;
s_mem_contents[14'h253e] = 8'h00;
s_mem_contents[14'h253f] = 8'h48;
s_mem_contents[14'h2540] = 8'hb5;
s_mem_contents[14'h2541] = 8'h09;
s_mem_contents[14'h2542] = 8'h8d;
s_mem_contents[14'h2543] = 8'h03;
s_mem_contents[14'h2544] = 8'h02;
s_mem_contents[14'h2545] = 8'h28;
s_mem_contents[14'h2546] = 8'h0e;
s_mem_contents[14'h2547] = 8'h03;
s_mem_contents[14'h2548] = 8'h02;
s_mem_contents[14'h2549] = 8'h08;
s_mem_contents[14'h254a] = 8'had;
s_mem_contents[14'h254b] = 8'h03;
s_mem_contents[14'h254c] = 8'h02;
s_mem_contents[14'h254d] = 8'hdd;
s_mem_contents[14'h254e] = 8'h20;
s_mem_contents[14'h254f] = 8'h02;
s_mem_contents[14'h2550] = 8'hd0;
s_mem_contents[14'h2551] = 8'hfe;
s_mem_contents[14'h2552] = 8'h68;
s_mem_contents[14'h2553] = 8'h49;
s_mem_contents[14'h2554] = 8'h30;
s_mem_contents[14'h2555] = 8'hdd;
s_mem_contents[14'h2556] = 8'h30;
s_mem_contents[14'h2557] = 8'h02;
s_mem_contents[14'h2558] = 8'hd0;
s_mem_contents[14'h2559] = 8'hfe;
s_mem_contents[14'h255a] = 8'hca;
s_mem_contents[14'h255b] = 8'h10;
s_mem_contents[14'h255c] = 8'he0;
s_mem_contents[14'h255d] = 8'ha2;
s_mem_contents[14'h255e] = 8'h03;
s_mem_contents[14'h255f] = 8'ha9;
s_mem_contents[14'h2560] = 8'hff;
s_mem_contents[14'h2561] = 8'h48;
s_mem_contents[14'h2562] = 8'hb5;
s_mem_contents[14'h2563] = 8'h09;
s_mem_contents[14'h2564] = 8'h8d;
s_mem_contents[14'h2565] = 8'h03;
s_mem_contents[14'h2566] = 8'h02;
s_mem_contents[14'h2567] = 8'h28;
s_mem_contents[14'h2568] = 8'h0e;
s_mem_contents[14'h2569] = 8'h03;
s_mem_contents[14'h256a] = 8'h02;
s_mem_contents[14'h256b] = 8'h08;
s_mem_contents[14'h256c] = 8'had;
s_mem_contents[14'h256d] = 8'h03;
s_mem_contents[14'h256e] = 8'h02;
s_mem_contents[14'h256f] = 8'hdd;
s_mem_contents[14'h2570] = 8'h20;
s_mem_contents[14'h2571] = 8'h02;
s_mem_contents[14'h2572] = 8'hd0;
s_mem_contents[14'h2573] = 8'hfe;
s_mem_contents[14'h2574] = 8'h68;
s_mem_contents[14'h2575] = 8'h49;
s_mem_contents[14'h2576] = 8'h7c;
s_mem_contents[14'h2577] = 8'hdd;
s_mem_contents[14'h2578] = 8'h30;
s_mem_contents[14'h2579] = 8'h02;
s_mem_contents[14'h257a] = 8'hd0;
s_mem_contents[14'h257b] = 8'hfe;
s_mem_contents[14'h257c] = 8'hca;
s_mem_contents[14'h257d] = 8'h10;
s_mem_contents[14'h257e] = 8'he0;
s_mem_contents[14'h257f] = 8'ha2;
s_mem_contents[14'h2580] = 8'h03;
s_mem_contents[14'h2581] = 8'ha9;
s_mem_contents[14'h2582] = 8'h00;
s_mem_contents[14'h2583] = 8'h48;
s_mem_contents[14'h2584] = 8'hb5;
s_mem_contents[14'h2585] = 8'h09;
s_mem_contents[14'h2586] = 8'h8d;
s_mem_contents[14'h2587] = 8'h03;
s_mem_contents[14'h2588] = 8'h02;
s_mem_contents[14'h2589] = 8'h28;
s_mem_contents[14'h258a] = 8'h4e;
s_mem_contents[14'h258b] = 8'h03;
s_mem_contents[14'h258c] = 8'h02;
s_mem_contents[14'h258d] = 8'h08;
s_mem_contents[14'h258e] = 8'had;
s_mem_contents[14'h258f] = 8'h03;
s_mem_contents[14'h2590] = 8'h02;
s_mem_contents[14'h2591] = 8'hdd;
s_mem_contents[14'h2592] = 8'h28;
s_mem_contents[14'h2593] = 8'h02;
s_mem_contents[14'h2594] = 8'hd0;
s_mem_contents[14'h2595] = 8'hfe;
s_mem_contents[14'h2596] = 8'h68;
s_mem_contents[14'h2597] = 8'h49;
s_mem_contents[14'h2598] = 8'h30;
s_mem_contents[14'h2599] = 8'hdd;
s_mem_contents[14'h259a] = 8'h38;
s_mem_contents[14'h259b] = 8'h02;
s_mem_contents[14'h259c] = 8'hd0;
s_mem_contents[14'h259d] = 8'hfe;
s_mem_contents[14'h259e] = 8'hca;
s_mem_contents[14'h259f] = 8'h10;
s_mem_contents[14'h25a0] = 8'he0;
s_mem_contents[14'h25a1] = 8'ha2;
s_mem_contents[14'h25a2] = 8'h03;
s_mem_contents[14'h25a3] = 8'ha9;
s_mem_contents[14'h25a4] = 8'hff;
s_mem_contents[14'h25a5] = 8'h48;
s_mem_contents[14'h25a6] = 8'hb5;
s_mem_contents[14'h25a7] = 8'h09;
s_mem_contents[14'h25a8] = 8'h8d;
s_mem_contents[14'h25a9] = 8'h03;
s_mem_contents[14'h25aa] = 8'h02;
s_mem_contents[14'h25ab] = 8'h28;
s_mem_contents[14'h25ac] = 8'h4e;
s_mem_contents[14'h25ad] = 8'h03;
s_mem_contents[14'h25ae] = 8'h02;
s_mem_contents[14'h25af] = 8'h08;
s_mem_contents[14'h25b0] = 8'had;
s_mem_contents[14'h25b1] = 8'h03;
s_mem_contents[14'h25b2] = 8'h02;
s_mem_contents[14'h25b3] = 8'hdd;
s_mem_contents[14'h25b4] = 8'h28;
s_mem_contents[14'h25b5] = 8'h02;
s_mem_contents[14'h25b6] = 8'hd0;
s_mem_contents[14'h25b7] = 8'hfe;
s_mem_contents[14'h25b8] = 8'h68;
s_mem_contents[14'h25b9] = 8'h49;
s_mem_contents[14'h25ba] = 8'h7c;
s_mem_contents[14'h25bb] = 8'hdd;
s_mem_contents[14'h25bc] = 8'h38;
s_mem_contents[14'h25bd] = 8'h02;
s_mem_contents[14'h25be] = 8'hd0;
s_mem_contents[14'h25bf] = 8'hfe;
s_mem_contents[14'h25c0] = 8'hca;
s_mem_contents[14'h25c1] = 8'h10;
s_mem_contents[14'h25c2] = 8'he0;
s_mem_contents[14'h25c3] = 8'ha2;
s_mem_contents[14'h25c4] = 8'h03;
s_mem_contents[14'h25c5] = 8'ha9;
s_mem_contents[14'h25c6] = 8'h00;
s_mem_contents[14'h25c7] = 8'h48;
s_mem_contents[14'h25c8] = 8'hb5;
s_mem_contents[14'h25c9] = 8'h09;
s_mem_contents[14'h25ca] = 8'h8d;
s_mem_contents[14'h25cb] = 8'h03;
s_mem_contents[14'h25cc] = 8'h02;
s_mem_contents[14'h25cd] = 8'h28;
s_mem_contents[14'h25ce] = 8'h2e;
s_mem_contents[14'h25cf] = 8'h03;
s_mem_contents[14'h25d0] = 8'h02;
s_mem_contents[14'h25d1] = 8'h08;
s_mem_contents[14'h25d2] = 8'had;
s_mem_contents[14'h25d3] = 8'h03;
s_mem_contents[14'h25d4] = 8'h02;
s_mem_contents[14'h25d5] = 8'hdd;
s_mem_contents[14'h25d6] = 8'h20;
s_mem_contents[14'h25d7] = 8'h02;
s_mem_contents[14'h25d8] = 8'hd0;
s_mem_contents[14'h25d9] = 8'hfe;
s_mem_contents[14'h25da] = 8'h68;
s_mem_contents[14'h25db] = 8'h49;
s_mem_contents[14'h25dc] = 8'h30;
s_mem_contents[14'h25dd] = 8'hdd;
s_mem_contents[14'h25de] = 8'h30;
s_mem_contents[14'h25df] = 8'h02;
s_mem_contents[14'h25e0] = 8'hd0;
s_mem_contents[14'h25e1] = 8'hfe;
s_mem_contents[14'h25e2] = 8'hca;
s_mem_contents[14'h25e3] = 8'h10;
s_mem_contents[14'h25e4] = 8'he0;
s_mem_contents[14'h25e5] = 8'ha2;
s_mem_contents[14'h25e6] = 8'h03;
s_mem_contents[14'h25e7] = 8'ha9;
s_mem_contents[14'h25e8] = 8'hfe;
s_mem_contents[14'h25e9] = 8'h48;
s_mem_contents[14'h25ea] = 8'hb5;
s_mem_contents[14'h25eb] = 8'h09;
s_mem_contents[14'h25ec] = 8'h8d;
s_mem_contents[14'h25ed] = 8'h03;
s_mem_contents[14'h25ee] = 8'h02;
s_mem_contents[14'h25ef] = 8'h28;
s_mem_contents[14'h25f0] = 8'h2e;
s_mem_contents[14'h25f1] = 8'h03;
s_mem_contents[14'h25f2] = 8'h02;
s_mem_contents[14'h25f3] = 8'h08;
s_mem_contents[14'h25f4] = 8'had;
s_mem_contents[14'h25f5] = 8'h03;
s_mem_contents[14'h25f6] = 8'h02;
s_mem_contents[14'h25f7] = 8'hdd;
s_mem_contents[14'h25f8] = 8'h20;
s_mem_contents[14'h25f9] = 8'h02;
s_mem_contents[14'h25fa] = 8'hd0;
s_mem_contents[14'h25fb] = 8'hfe;
s_mem_contents[14'h25fc] = 8'h68;
s_mem_contents[14'h25fd] = 8'h49;
s_mem_contents[14'h25fe] = 8'h7c;
s_mem_contents[14'h25ff] = 8'hdd;
s_mem_contents[14'h2600] = 8'h30;
s_mem_contents[14'h2601] = 8'h02;
s_mem_contents[14'h2602] = 8'hd0;
s_mem_contents[14'h2603] = 8'hfe;
s_mem_contents[14'h2604] = 8'hca;
s_mem_contents[14'h2605] = 8'h10;
s_mem_contents[14'h2606] = 8'he0;
s_mem_contents[14'h2607] = 8'ha2;
s_mem_contents[14'h2608] = 8'h03;
s_mem_contents[14'h2609] = 8'ha9;
s_mem_contents[14'h260a] = 8'h01;
s_mem_contents[14'h260b] = 8'h48;
s_mem_contents[14'h260c] = 8'hb5;
s_mem_contents[14'h260d] = 8'h09;
s_mem_contents[14'h260e] = 8'h8d;
s_mem_contents[14'h260f] = 8'h03;
s_mem_contents[14'h2610] = 8'h02;
s_mem_contents[14'h2611] = 8'h28;
s_mem_contents[14'h2612] = 8'h2e;
s_mem_contents[14'h2613] = 8'h03;
s_mem_contents[14'h2614] = 8'h02;
s_mem_contents[14'h2615] = 8'h08;
s_mem_contents[14'h2616] = 8'had;
s_mem_contents[14'h2617] = 8'h03;
s_mem_contents[14'h2618] = 8'h02;
s_mem_contents[14'h2619] = 8'hdd;
s_mem_contents[14'h261a] = 8'h24;
s_mem_contents[14'h261b] = 8'h02;
s_mem_contents[14'h261c] = 8'hd0;
s_mem_contents[14'h261d] = 8'hfe;
s_mem_contents[14'h261e] = 8'h68;
s_mem_contents[14'h261f] = 8'h49;
s_mem_contents[14'h2620] = 8'h30;
s_mem_contents[14'h2621] = 8'hdd;
s_mem_contents[14'h2622] = 8'h34;
s_mem_contents[14'h2623] = 8'h02;
s_mem_contents[14'h2624] = 8'hd0;
s_mem_contents[14'h2625] = 8'hfe;
s_mem_contents[14'h2626] = 8'hca;
s_mem_contents[14'h2627] = 8'h10;
s_mem_contents[14'h2628] = 8'he0;
s_mem_contents[14'h2629] = 8'ha2;
s_mem_contents[14'h262a] = 8'h03;
s_mem_contents[14'h262b] = 8'ha9;
s_mem_contents[14'h262c] = 8'hff;
s_mem_contents[14'h262d] = 8'h48;
s_mem_contents[14'h262e] = 8'hb5;
s_mem_contents[14'h262f] = 8'h09;
s_mem_contents[14'h2630] = 8'h8d;
s_mem_contents[14'h2631] = 8'h03;
s_mem_contents[14'h2632] = 8'h02;
s_mem_contents[14'h2633] = 8'h28;
s_mem_contents[14'h2634] = 8'h2e;
s_mem_contents[14'h2635] = 8'h03;
s_mem_contents[14'h2636] = 8'h02;
s_mem_contents[14'h2637] = 8'h08;
s_mem_contents[14'h2638] = 8'had;
s_mem_contents[14'h2639] = 8'h03;
s_mem_contents[14'h263a] = 8'h02;
s_mem_contents[14'h263b] = 8'hdd;
s_mem_contents[14'h263c] = 8'h24;
s_mem_contents[14'h263d] = 8'h02;
s_mem_contents[14'h263e] = 8'hd0;
s_mem_contents[14'h263f] = 8'hfe;
s_mem_contents[14'h2640] = 8'h68;
s_mem_contents[14'h2641] = 8'h49;
s_mem_contents[14'h2642] = 8'h7c;
s_mem_contents[14'h2643] = 8'hdd;
s_mem_contents[14'h2644] = 8'h34;
s_mem_contents[14'h2645] = 8'h02;
s_mem_contents[14'h2646] = 8'hd0;
s_mem_contents[14'h2647] = 8'hfe;
s_mem_contents[14'h2648] = 8'hca;
s_mem_contents[14'h2649] = 8'h10;
s_mem_contents[14'h264a] = 8'he0;
s_mem_contents[14'h264b] = 8'ha2;
s_mem_contents[14'h264c] = 8'h03;
s_mem_contents[14'h264d] = 8'ha9;
s_mem_contents[14'h264e] = 8'h00;
s_mem_contents[14'h264f] = 8'h48;
s_mem_contents[14'h2650] = 8'hb5;
s_mem_contents[14'h2651] = 8'h09;
s_mem_contents[14'h2652] = 8'h8d;
s_mem_contents[14'h2653] = 8'h03;
s_mem_contents[14'h2654] = 8'h02;
s_mem_contents[14'h2655] = 8'h28;
s_mem_contents[14'h2656] = 8'h6e;
s_mem_contents[14'h2657] = 8'h03;
s_mem_contents[14'h2658] = 8'h02;
s_mem_contents[14'h2659] = 8'h08;
s_mem_contents[14'h265a] = 8'had;
s_mem_contents[14'h265b] = 8'h03;
s_mem_contents[14'h265c] = 8'h02;
s_mem_contents[14'h265d] = 8'hdd;
s_mem_contents[14'h265e] = 8'h28;
s_mem_contents[14'h265f] = 8'h02;
s_mem_contents[14'h2660] = 8'hd0;
s_mem_contents[14'h2661] = 8'hfe;
s_mem_contents[14'h2662] = 8'h68;
s_mem_contents[14'h2663] = 8'h49;
s_mem_contents[14'h2664] = 8'h30;
s_mem_contents[14'h2665] = 8'hdd;
s_mem_contents[14'h2666] = 8'h38;
s_mem_contents[14'h2667] = 8'h02;
s_mem_contents[14'h2668] = 8'hd0;
s_mem_contents[14'h2669] = 8'hfe;
s_mem_contents[14'h266a] = 8'hca;
s_mem_contents[14'h266b] = 8'h10;
s_mem_contents[14'h266c] = 8'he0;
s_mem_contents[14'h266d] = 8'ha2;
s_mem_contents[14'h266e] = 8'h03;
s_mem_contents[14'h266f] = 8'ha9;
s_mem_contents[14'h2670] = 8'hfe;
s_mem_contents[14'h2671] = 8'h48;
s_mem_contents[14'h2672] = 8'hb5;
s_mem_contents[14'h2673] = 8'h09;
s_mem_contents[14'h2674] = 8'h8d;
s_mem_contents[14'h2675] = 8'h03;
s_mem_contents[14'h2676] = 8'h02;
s_mem_contents[14'h2677] = 8'h28;
s_mem_contents[14'h2678] = 8'h6e;
s_mem_contents[14'h2679] = 8'h03;
s_mem_contents[14'h267a] = 8'h02;
s_mem_contents[14'h267b] = 8'h08;
s_mem_contents[14'h267c] = 8'had;
s_mem_contents[14'h267d] = 8'h03;
s_mem_contents[14'h267e] = 8'h02;
s_mem_contents[14'h267f] = 8'hdd;
s_mem_contents[14'h2680] = 8'h28;
s_mem_contents[14'h2681] = 8'h02;
s_mem_contents[14'h2682] = 8'hd0;
s_mem_contents[14'h2683] = 8'hfe;
s_mem_contents[14'h2684] = 8'h68;
s_mem_contents[14'h2685] = 8'h49;
s_mem_contents[14'h2686] = 8'h7c;
s_mem_contents[14'h2687] = 8'hdd;
s_mem_contents[14'h2688] = 8'h38;
s_mem_contents[14'h2689] = 8'h02;
s_mem_contents[14'h268a] = 8'hd0;
s_mem_contents[14'h268b] = 8'hfe;
s_mem_contents[14'h268c] = 8'hca;
s_mem_contents[14'h268d] = 8'h10;
s_mem_contents[14'h268e] = 8'he0;
s_mem_contents[14'h268f] = 8'ha2;
s_mem_contents[14'h2690] = 8'h03;
s_mem_contents[14'h2691] = 8'ha9;
s_mem_contents[14'h2692] = 8'h01;
s_mem_contents[14'h2693] = 8'h48;
s_mem_contents[14'h2694] = 8'hb5;
s_mem_contents[14'h2695] = 8'h09;
s_mem_contents[14'h2696] = 8'h8d;
s_mem_contents[14'h2697] = 8'h03;
s_mem_contents[14'h2698] = 8'h02;
s_mem_contents[14'h2699] = 8'h28;
s_mem_contents[14'h269a] = 8'h6e;
s_mem_contents[14'h269b] = 8'h03;
s_mem_contents[14'h269c] = 8'h02;
s_mem_contents[14'h269d] = 8'h08;
s_mem_contents[14'h269e] = 8'had;
s_mem_contents[14'h269f] = 8'h03;
s_mem_contents[14'h26a0] = 8'h02;
s_mem_contents[14'h26a1] = 8'hdd;
s_mem_contents[14'h26a2] = 8'h2c;
s_mem_contents[14'h26a3] = 8'h02;
s_mem_contents[14'h26a4] = 8'hd0;
s_mem_contents[14'h26a5] = 8'hfe;
s_mem_contents[14'h26a6] = 8'h68;
s_mem_contents[14'h26a7] = 8'h49;
s_mem_contents[14'h26a8] = 8'h30;
s_mem_contents[14'h26a9] = 8'hdd;
s_mem_contents[14'h26aa] = 8'h3c;
s_mem_contents[14'h26ab] = 8'h02;
s_mem_contents[14'h26ac] = 8'hd0;
s_mem_contents[14'h26ad] = 8'hfe;
s_mem_contents[14'h26ae] = 8'hca;
s_mem_contents[14'h26af] = 8'h10;
s_mem_contents[14'h26b0] = 8'he0;
s_mem_contents[14'h26b1] = 8'ha2;
s_mem_contents[14'h26b2] = 8'h03;
s_mem_contents[14'h26b3] = 8'ha9;
s_mem_contents[14'h26b4] = 8'hff;
s_mem_contents[14'h26b5] = 8'h48;
s_mem_contents[14'h26b6] = 8'hb5;
s_mem_contents[14'h26b7] = 8'h09;
s_mem_contents[14'h26b8] = 8'h8d;
s_mem_contents[14'h26b9] = 8'h03;
s_mem_contents[14'h26ba] = 8'h02;
s_mem_contents[14'h26bb] = 8'h28;
s_mem_contents[14'h26bc] = 8'h6e;
s_mem_contents[14'h26bd] = 8'h03;
s_mem_contents[14'h26be] = 8'h02;
s_mem_contents[14'h26bf] = 8'h08;
s_mem_contents[14'h26c0] = 8'had;
s_mem_contents[14'h26c1] = 8'h03;
s_mem_contents[14'h26c2] = 8'h02;
s_mem_contents[14'h26c3] = 8'hdd;
s_mem_contents[14'h26c4] = 8'h2c;
s_mem_contents[14'h26c5] = 8'h02;
s_mem_contents[14'h26c6] = 8'hd0;
s_mem_contents[14'h26c7] = 8'hfe;
s_mem_contents[14'h26c8] = 8'h68;
s_mem_contents[14'h26c9] = 8'h49;
s_mem_contents[14'h26ca] = 8'h7c;
s_mem_contents[14'h26cb] = 8'hdd;
s_mem_contents[14'h26cc] = 8'h3c;
s_mem_contents[14'h26cd] = 8'h02;
s_mem_contents[14'h26ce] = 8'hd0;
s_mem_contents[14'h26cf] = 8'hfe;
s_mem_contents[14'h26d0] = 8'hca;
s_mem_contents[14'h26d1] = 8'h10;
s_mem_contents[14'h26d2] = 8'he0;
s_mem_contents[14'h26d3] = 8'had;
s_mem_contents[14'h26d4] = 8'h00;
s_mem_contents[14'h26d5] = 8'h02;
s_mem_contents[14'h26d6] = 8'hc9;
s_mem_contents[14'h26d7] = 8'h1f;
s_mem_contents[14'h26d8] = 8'hd0;
s_mem_contents[14'h26d9] = 8'hfe;
s_mem_contents[14'h26da] = 8'ha9;
s_mem_contents[14'h26db] = 8'h20;
s_mem_contents[14'h26dc] = 8'h8d;
s_mem_contents[14'h26dd] = 8'h00;
s_mem_contents[14'h26de] = 8'h02;
s_mem_contents[14'h26df] = 8'ha2;
s_mem_contents[14'h26e0] = 8'h03;
s_mem_contents[14'h26e1] = 8'ha9;
s_mem_contents[14'h26e2] = 8'h00;
s_mem_contents[14'h26e3] = 8'h48;
s_mem_contents[14'h26e4] = 8'hb5;
s_mem_contents[14'h26e5] = 8'h09;
s_mem_contents[14'h26e6] = 8'h95;
s_mem_contents[14'h26e7] = 8'h02;
s_mem_contents[14'h26e8] = 8'h28;
s_mem_contents[14'h26e9] = 8'h16;
s_mem_contents[14'h26ea] = 8'h02;
s_mem_contents[14'h26eb] = 8'h08;
s_mem_contents[14'h26ec] = 8'hb5;
s_mem_contents[14'h26ed] = 8'h02;
s_mem_contents[14'h26ee] = 8'hdd;
s_mem_contents[14'h26ef] = 8'h20;
s_mem_contents[14'h26f0] = 8'h02;
s_mem_contents[14'h26f1] = 8'hd0;
s_mem_contents[14'h26f2] = 8'hfe;
s_mem_contents[14'h26f3] = 8'h68;
s_mem_contents[14'h26f4] = 8'h49;
s_mem_contents[14'h26f5] = 8'h30;
s_mem_contents[14'h26f6] = 8'hdd;
s_mem_contents[14'h26f7] = 8'h30;
s_mem_contents[14'h26f8] = 8'h02;
s_mem_contents[14'h26f9] = 8'hd0;
s_mem_contents[14'h26fa] = 8'hfe;
s_mem_contents[14'h26fb] = 8'hca;
s_mem_contents[14'h26fc] = 8'h10;
s_mem_contents[14'h26fd] = 8'he3;
s_mem_contents[14'h26fe] = 8'ha2;
s_mem_contents[14'h26ff] = 8'h03;
s_mem_contents[14'h2700] = 8'ha9;
s_mem_contents[14'h2701] = 8'hff;
s_mem_contents[14'h2702] = 8'h48;
s_mem_contents[14'h2703] = 8'hb5;
s_mem_contents[14'h2704] = 8'h09;
s_mem_contents[14'h2705] = 8'h95;
s_mem_contents[14'h2706] = 8'h02;
s_mem_contents[14'h2707] = 8'h28;
s_mem_contents[14'h2708] = 8'h16;
s_mem_contents[14'h2709] = 8'h02;
s_mem_contents[14'h270a] = 8'h08;
s_mem_contents[14'h270b] = 8'hb5;
s_mem_contents[14'h270c] = 8'h02;
s_mem_contents[14'h270d] = 8'hdd;
s_mem_contents[14'h270e] = 8'h20;
s_mem_contents[14'h270f] = 8'h02;
s_mem_contents[14'h2710] = 8'hd0;
s_mem_contents[14'h2711] = 8'hfe;
s_mem_contents[14'h2712] = 8'h68;
s_mem_contents[14'h2713] = 8'h49;
s_mem_contents[14'h2714] = 8'h7c;
s_mem_contents[14'h2715] = 8'hdd;
s_mem_contents[14'h2716] = 8'h30;
s_mem_contents[14'h2717] = 8'h02;
s_mem_contents[14'h2718] = 8'hd0;
s_mem_contents[14'h2719] = 8'hfe;
s_mem_contents[14'h271a] = 8'hca;
s_mem_contents[14'h271b] = 8'h10;
s_mem_contents[14'h271c] = 8'he3;
s_mem_contents[14'h271d] = 8'ha2;
s_mem_contents[14'h271e] = 8'h03;
s_mem_contents[14'h271f] = 8'ha9;
s_mem_contents[14'h2720] = 8'h00;
s_mem_contents[14'h2721] = 8'h48;
s_mem_contents[14'h2722] = 8'hb5;
s_mem_contents[14'h2723] = 8'h09;
s_mem_contents[14'h2724] = 8'h95;
s_mem_contents[14'h2725] = 8'h02;
s_mem_contents[14'h2726] = 8'h28;
s_mem_contents[14'h2727] = 8'h56;
s_mem_contents[14'h2728] = 8'h02;
s_mem_contents[14'h2729] = 8'h08;
s_mem_contents[14'h272a] = 8'hb5;
s_mem_contents[14'h272b] = 8'h02;
s_mem_contents[14'h272c] = 8'hdd;
s_mem_contents[14'h272d] = 8'h28;
s_mem_contents[14'h272e] = 8'h02;
s_mem_contents[14'h272f] = 8'hd0;
s_mem_contents[14'h2730] = 8'hfe;
s_mem_contents[14'h2731] = 8'h68;
s_mem_contents[14'h2732] = 8'h49;
s_mem_contents[14'h2733] = 8'h30;
s_mem_contents[14'h2734] = 8'hdd;
s_mem_contents[14'h2735] = 8'h38;
s_mem_contents[14'h2736] = 8'h02;
s_mem_contents[14'h2737] = 8'hd0;
s_mem_contents[14'h2738] = 8'hfe;
s_mem_contents[14'h2739] = 8'hca;
s_mem_contents[14'h273a] = 8'h10;
s_mem_contents[14'h273b] = 8'he3;
s_mem_contents[14'h273c] = 8'ha2;
s_mem_contents[14'h273d] = 8'h03;
s_mem_contents[14'h273e] = 8'ha9;
s_mem_contents[14'h273f] = 8'hff;
s_mem_contents[14'h2740] = 8'h48;
s_mem_contents[14'h2741] = 8'hb5;
s_mem_contents[14'h2742] = 8'h09;
s_mem_contents[14'h2743] = 8'h95;
s_mem_contents[14'h2744] = 8'h02;
s_mem_contents[14'h2745] = 8'h28;
s_mem_contents[14'h2746] = 8'h56;
s_mem_contents[14'h2747] = 8'h02;
s_mem_contents[14'h2748] = 8'h08;
s_mem_contents[14'h2749] = 8'hb5;
s_mem_contents[14'h274a] = 8'h02;
s_mem_contents[14'h274b] = 8'hdd;
s_mem_contents[14'h274c] = 8'h28;
s_mem_contents[14'h274d] = 8'h02;
s_mem_contents[14'h274e] = 8'hd0;
s_mem_contents[14'h274f] = 8'hfe;
s_mem_contents[14'h2750] = 8'h68;
s_mem_contents[14'h2751] = 8'h49;
s_mem_contents[14'h2752] = 8'h7c;
s_mem_contents[14'h2753] = 8'hdd;
s_mem_contents[14'h2754] = 8'h38;
s_mem_contents[14'h2755] = 8'h02;
s_mem_contents[14'h2756] = 8'hd0;
s_mem_contents[14'h2757] = 8'hfe;
s_mem_contents[14'h2758] = 8'hca;
s_mem_contents[14'h2759] = 8'h10;
s_mem_contents[14'h275a] = 8'he3;
s_mem_contents[14'h275b] = 8'ha2;
s_mem_contents[14'h275c] = 8'h03;
s_mem_contents[14'h275d] = 8'ha9;
s_mem_contents[14'h275e] = 8'h00;
s_mem_contents[14'h275f] = 8'h48;
s_mem_contents[14'h2760] = 8'hb5;
s_mem_contents[14'h2761] = 8'h09;
s_mem_contents[14'h2762] = 8'h95;
s_mem_contents[14'h2763] = 8'h02;
s_mem_contents[14'h2764] = 8'h28;
s_mem_contents[14'h2765] = 8'h36;
s_mem_contents[14'h2766] = 8'h02;
s_mem_contents[14'h2767] = 8'h08;
s_mem_contents[14'h2768] = 8'hb5;
s_mem_contents[14'h2769] = 8'h02;
s_mem_contents[14'h276a] = 8'hdd;
s_mem_contents[14'h276b] = 8'h20;
s_mem_contents[14'h276c] = 8'h02;
s_mem_contents[14'h276d] = 8'hd0;
s_mem_contents[14'h276e] = 8'hfe;
s_mem_contents[14'h276f] = 8'h68;
s_mem_contents[14'h2770] = 8'h49;
s_mem_contents[14'h2771] = 8'h30;
s_mem_contents[14'h2772] = 8'hdd;
s_mem_contents[14'h2773] = 8'h30;
s_mem_contents[14'h2774] = 8'h02;
s_mem_contents[14'h2775] = 8'hd0;
s_mem_contents[14'h2776] = 8'hfe;
s_mem_contents[14'h2777] = 8'hca;
s_mem_contents[14'h2778] = 8'h10;
s_mem_contents[14'h2779] = 8'he3;
s_mem_contents[14'h277a] = 8'ha2;
s_mem_contents[14'h277b] = 8'h03;
s_mem_contents[14'h277c] = 8'ha9;
s_mem_contents[14'h277d] = 8'hfe;
s_mem_contents[14'h277e] = 8'h48;
s_mem_contents[14'h277f] = 8'hb5;
s_mem_contents[14'h2780] = 8'h09;
s_mem_contents[14'h2781] = 8'h95;
s_mem_contents[14'h2782] = 8'h02;
s_mem_contents[14'h2783] = 8'h28;
s_mem_contents[14'h2784] = 8'h36;
s_mem_contents[14'h2785] = 8'h02;
s_mem_contents[14'h2786] = 8'h08;
s_mem_contents[14'h2787] = 8'hb5;
s_mem_contents[14'h2788] = 8'h02;
s_mem_contents[14'h2789] = 8'hdd;
s_mem_contents[14'h278a] = 8'h20;
s_mem_contents[14'h278b] = 8'h02;
s_mem_contents[14'h278c] = 8'hd0;
s_mem_contents[14'h278d] = 8'hfe;
s_mem_contents[14'h278e] = 8'h68;
s_mem_contents[14'h278f] = 8'h49;
s_mem_contents[14'h2790] = 8'h7c;
s_mem_contents[14'h2791] = 8'hdd;
s_mem_contents[14'h2792] = 8'h30;
s_mem_contents[14'h2793] = 8'h02;
s_mem_contents[14'h2794] = 8'hd0;
s_mem_contents[14'h2795] = 8'hfe;
s_mem_contents[14'h2796] = 8'hca;
s_mem_contents[14'h2797] = 8'h10;
s_mem_contents[14'h2798] = 8'he3;
s_mem_contents[14'h2799] = 8'ha2;
s_mem_contents[14'h279a] = 8'h03;
s_mem_contents[14'h279b] = 8'ha9;
s_mem_contents[14'h279c] = 8'h01;
s_mem_contents[14'h279d] = 8'h48;
s_mem_contents[14'h279e] = 8'hb5;
s_mem_contents[14'h279f] = 8'h09;
s_mem_contents[14'h27a0] = 8'h95;
s_mem_contents[14'h27a1] = 8'h02;
s_mem_contents[14'h27a2] = 8'h28;
s_mem_contents[14'h27a3] = 8'h36;
s_mem_contents[14'h27a4] = 8'h02;
s_mem_contents[14'h27a5] = 8'h08;
s_mem_contents[14'h27a6] = 8'hb5;
s_mem_contents[14'h27a7] = 8'h02;
s_mem_contents[14'h27a8] = 8'hdd;
s_mem_contents[14'h27a9] = 8'h24;
s_mem_contents[14'h27aa] = 8'h02;
s_mem_contents[14'h27ab] = 8'hd0;
s_mem_contents[14'h27ac] = 8'hfe;
s_mem_contents[14'h27ad] = 8'h68;
s_mem_contents[14'h27ae] = 8'h49;
s_mem_contents[14'h27af] = 8'h30;
s_mem_contents[14'h27b0] = 8'hdd;
s_mem_contents[14'h27b1] = 8'h34;
s_mem_contents[14'h27b2] = 8'h02;
s_mem_contents[14'h27b3] = 8'hd0;
s_mem_contents[14'h27b4] = 8'hfe;
s_mem_contents[14'h27b5] = 8'hca;
s_mem_contents[14'h27b6] = 8'h10;
s_mem_contents[14'h27b7] = 8'he3;
s_mem_contents[14'h27b8] = 8'ha2;
s_mem_contents[14'h27b9] = 8'h03;
s_mem_contents[14'h27ba] = 8'ha9;
s_mem_contents[14'h27bb] = 8'hff;
s_mem_contents[14'h27bc] = 8'h48;
s_mem_contents[14'h27bd] = 8'hb5;
s_mem_contents[14'h27be] = 8'h09;
s_mem_contents[14'h27bf] = 8'h95;
s_mem_contents[14'h27c0] = 8'h02;
s_mem_contents[14'h27c1] = 8'h28;
s_mem_contents[14'h27c2] = 8'h36;
s_mem_contents[14'h27c3] = 8'h02;
s_mem_contents[14'h27c4] = 8'h08;
s_mem_contents[14'h27c5] = 8'hb5;
s_mem_contents[14'h27c6] = 8'h02;
s_mem_contents[14'h27c7] = 8'hdd;
s_mem_contents[14'h27c8] = 8'h24;
s_mem_contents[14'h27c9] = 8'h02;
s_mem_contents[14'h27ca] = 8'hd0;
s_mem_contents[14'h27cb] = 8'hfe;
s_mem_contents[14'h27cc] = 8'h68;
s_mem_contents[14'h27cd] = 8'h49;
s_mem_contents[14'h27ce] = 8'h7c;
s_mem_contents[14'h27cf] = 8'hdd;
s_mem_contents[14'h27d0] = 8'h34;
s_mem_contents[14'h27d1] = 8'h02;
s_mem_contents[14'h27d2] = 8'hd0;
s_mem_contents[14'h27d3] = 8'hfe;
s_mem_contents[14'h27d4] = 8'hca;
s_mem_contents[14'h27d5] = 8'h10;
s_mem_contents[14'h27d6] = 8'he3;
s_mem_contents[14'h27d7] = 8'ha2;
s_mem_contents[14'h27d8] = 8'h03;
s_mem_contents[14'h27d9] = 8'ha9;
s_mem_contents[14'h27da] = 8'h00;
s_mem_contents[14'h27db] = 8'h48;
s_mem_contents[14'h27dc] = 8'hb5;
s_mem_contents[14'h27dd] = 8'h09;
s_mem_contents[14'h27de] = 8'h95;
s_mem_contents[14'h27df] = 8'h02;
s_mem_contents[14'h27e0] = 8'h28;
s_mem_contents[14'h27e1] = 8'h76;
s_mem_contents[14'h27e2] = 8'h02;
s_mem_contents[14'h27e3] = 8'h08;
s_mem_contents[14'h27e4] = 8'hb5;
s_mem_contents[14'h27e5] = 8'h02;
s_mem_contents[14'h27e6] = 8'hdd;
s_mem_contents[14'h27e7] = 8'h28;
s_mem_contents[14'h27e8] = 8'h02;
s_mem_contents[14'h27e9] = 8'hd0;
s_mem_contents[14'h27ea] = 8'hfe;
s_mem_contents[14'h27eb] = 8'h68;
s_mem_contents[14'h27ec] = 8'h49;
s_mem_contents[14'h27ed] = 8'h30;
s_mem_contents[14'h27ee] = 8'hdd;
s_mem_contents[14'h27ef] = 8'h38;
s_mem_contents[14'h27f0] = 8'h02;
s_mem_contents[14'h27f1] = 8'hd0;
s_mem_contents[14'h27f2] = 8'hfe;
s_mem_contents[14'h27f3] = 8'hca;
s_mem_contents[14'h27f4] = 8'h10;
s_mem_contents[14'h27f5] = 8'he3;
s_mem_contents[14'h27f6] = 8'ha2;
s_mem_contents[14'h27f7] = 8'h03;
s_mem_contents[14'h27f8] = 8'ha9;
s_mem_contents[14'h27f9] = 8'hfe;
s_mem_contents[14'h27fa] = 8'h48;
s_mem_contents[14'h27fb] = 8'hb5;
s_mem_contents[14'h27fc] = 8'h09;
s_mem_contents[14'h27fd] = 8'h95;
s_mem_contents[14'h27fe] = 8'h02;
s_mem_contents[14'h27ff] = 8'h28;
s_mem_contents[14'h2800] = 8'h76;
s_mem_contents[14'h2801] = 8'h02;
s_mem_contents[14'h2802] = 8'h08;
s_mem_contents[14'h2803] = 8'hb5;
s_mem_contents[14'h2804] = 8'h02;
s_mem_contents[14'h2805] = 8'hdd;
s_mem_contents[14'h2806] = 8'h28;
s_mem_contents[14'h2807] = 8'h02;
s_mem_contents[14'h2808] = 8'hd0;
s_mem_contents[14'h2809] = 8'hfe;
s_mem_contents[14'h280a] = 8'h68;
s_mem_contents[14'h280b] = 8'h49;
s_mem_contents[14'h280c] = 8'h7c;
s_mem_contents[14'h280d] = 8'hdd;
s_mem_contents[14'h280e] = 8'h38;
s_mem_contents[14'h280f] = 8'h02;
s_mem_contents[14'h2810] = 8'hd0;
s_mem_contents[14'h2811] = 8'hfe;
s_mem_contents[14'h2812] = 8'hca;
s_mem_contents[14'h2813] = 8'h10;
s_mem_contents[14'h2814] = 8'he3;
s_mem_contents[14'h2815] = 8'ha2;
s_mem_contents[14'h2816] = 8'h03;
s_mem_contents[14'h2817] = 8'ha9;
s_mem_contents[14'h2818] = 8'h01;
s_mem_contents[14'h2819] = 8'h48;
s_mem_contents[14'h281a] = 8'hb5;
s_mem_contents[14'h281b] = 8'h09;
s_mem_contents[14'h281c] = 8'h95;
s_mem_contents[14'h281d] = 8'h02;
s_mem_contents[14'h281e] = 8'h28;
s_mem_contents[14'h281f] = 8'h76;
s_mem_contents[14'h2820] = 8'h02;
s_mem_contents[14'h2821] = 8'h08;
s_mem_contents[14'h2822] = 8'hb5;
s_mem_contents[14'h2823] = 8'h02;
s_mem_contents[14'h2824] = 8'hdd;
s_mem_contents[14'h2825] = 8'h2c;
s_mem_contents[14'h2826] = 8'h02;
s_mem_contents[14'h2827] = 8'hd0;
s_mem_contents[14'h2828] = 8'hfe;
s_mem_contents[14'h2829] = 8'h68;
s_mem_contents[14'h282a] = 8'h49;
s_mem_contents[14'h282b] = 8'h30;
s_mem_contents[14'h282c] = 8'hdd;
s_mem_contents[14'h282d] = 8'h3c;
s_mem_contents[14'h282e] = 8'h02;
s_mem_contents[14'h282f] = 8'hd0;
s_mem_contents[14'h2830] = 8'hfe;
s_mem_contents[14'h2831] = 8'hca;
s_mem_contents[14'h2832] = 8'h10;
s_mem_contents[14'h2833] = 8'he3;
s_mem_contents[14'h2834] = 8'ha2;
s_mem_contents[14'h2835] = 8'h03;
s_mem_contents[14'h2836] = 8'ha9;
s_mem_contents[14'h2837] = 8'hff;
s_mem_contents[14'h2838] = 8'h48;
s_mem_contents[14'h2839] = 8'hb5;
s_mem_contents[14'h283a] = 8'h09;
s_mem_contents[14'h283b] = 8'h95;
s_mem_contents[14'h283c] = 8'h02;
s_mem_contents[14'h283d] = 8'h28;
s_mem_contents[14'h283e] = 8'h76;
s_mem_contents[14'h283f] = 8'h02;
s_mem_contents[14'h2840] = 8'h08;
s_mem_contents[14'h2841] = 8'hb5;
s_mem_contents[14'h2842] = 8'h02;
s_mem_contents[14'h2843] = 8'hdd;
s_mem_contents[14'h2844] = 8'h2c;
s_mem_contents[14'h2845] = 8'h02;
s_mem_contents[14'h2846] = 8'hd0;
s_mem_contents[14'h2847] = 8'hfe;
s_mem_contents[14'h2848] = 8'h68;
s_mem_contents[14'h2849] = 8'h49;
s_mem_contents[14'h284a] = 8'h7c;
s_mem_contents[14'h284b] = 8'hdd;
s_mem_contents[14'h284c] = 8'h3c;
s_mem_contents[14'h284d] = 8'h02;
s_mem_contents[14'h284e] = 8'hd0;
s_mem_contents[14'h284f] = 8'hfe;
s_mem_contents[14'h2850] = 8'hca;
s_mem_contents[14'h2851] = 8'h10;
s_mem_contents[14'h2852] = 8'he3;
s_mem_contents[14'h2853] = 8'had;
s_mem_contents[14'h2854] = 8'h00;
s_mem_contents[14'h2855] = 8'h02;
s_mem_contents[14'h2856] = 8'hc9;
s_mem_contents[14'h2857] = 8'h20;
s_mem_contents[14'h2858] = 8'hd0;
s_mem_contents[14'h2859] = 8'hfe;
s_mem_contents[14'h285a] = 8'ha9;
s_mem_contents[14'h285b] = 8'h21;
s_mem_contents[14'h285c] = 8'h8d;
s_mem_contents[14'h285d] = 8'h00;
s_mem_contents[14'h285e] = 8'h02;
s_mem_contents[14'h285f] = 8'ha2;
s_mem_contents[14'h2860] = 8'h03;
s_mem_contents[14'h2861] = 8'ha9;
s_mem_contents[14'h2862] = 8'h00;
s_mem_contents[14'h2863] = 8'h48;
s_mem_contents[14'h2864] = 8'hb5;
s_mem_contents[14'h2865] = 8'h09;
s_mem_contents[14'h2866] = 8'h9d;
s_mem_contents[14'h2867] = 8'h03;
s_mem_contents[14'h2868] = 8'h02;
s_mem_contents[14'h2869] = 8'h28;
s_mem_contents[14'h286a] = 8'h1e;
s_mem_contents[14'h286b] = 8'h03;
s_mem_contents[14'h286c] = 8'h02;
s_mem_contents[14'h286d] = 8'h08;
s_mem_contents[14'h286e] = 8'hbd;
s_mem_contents[14'h286f] = 8'h03;
s_mem_contents[14'h2870] = 8'h02;
s_mem_contents[14'h2871] = 8'hdd;
s_mem_contents[14'h2872] = 8'h20;
s_mem_contents[14'h2873] = 8'h02;
s_mem_contents[14'h2874] = 8'hd0;
s_mem_contents[14'h2875] = 8'hfe;
s_mem_contents[14'h2876] = 8'h68;
s_mem_contents[14'h2877] = 8'h49;
s_mem_contents[14'h2878] = 8'h30;
s_mem_contents[14'h2879] = 8'hdd;
s_mem_contents[14'h287a] = 8'h30;
s_mem_contents[14'h287b] = 8'h02;
s_mem_contents[14'h287c] = 8'hd0;
s_mem_contents[14'h287d] = 8'hfe;
s_mem_contents[14'h287e] = 8'hca;
s_mem_contents[14'h287f] = 8'h10;
s_mem_contents[14'h2880] = 8'he0;
s_mem_contents[14'h2881] = 8'ha2;
s_mem_contents[14'h2882] = 8'h03;
s_mem_contents[14'h2883] = 8'ha9;
s_mem_contents[14'h2884] = 8'hff;
s_mem_contents[14'h2885] = 8'h48;
s_mem_contents[14'h2886] = 8'hb5;
s_mem_contents[14'h2887] = 8'h09;
s_mem_contents[14'h2888] = 8'h9d;
s_mem_contents[14'h2889] = 8'h03;
s_mem_contents[14'h288a] = 8'h02;
s_mem_contents[14'h288b] = 8'h28;
s_mem_contents[14'h288c] = 8'h1e;
s_mem_contents[14'h288d] = 8'h03;
s_mem_contents[14'h288e] = 8'h02;
s_mem_contents[14'h288f] = 8'h08;
s_mem_contents[14'h2890] = 8'hbd;
s_mem_contents[14'h2891] = 8'h03;
s_mem_contents[14'h2892] = 8'h02;
s_mem_contents[14'h2893] = 8'hdd;
s_mem_contents[14'h2894] = 8'h20;
s_mem_contents[14'h2895] = 8'h02;
s_mem_contents[14'h2896] = 8'hd0;
s_mem_contents[14'h2897] = 8'hfe;
s_mem_contents[14'h2898] = 8'h68;
s_mem_contents[14'h2899] = 8'h49;
s_mem_contents[14'h289a] = 8'h7c;
s_mem_contents[14'h289b] = 8'hdd;
s_mem_contents[14'h289c] = 8'h30;
s_mem_contents[14'h289d] = 8'h02;
s_mem_contents[14'h289e] = 8'hd0;
s_mem_contents[14'h289f] = 8'hfe;
s_mem_contents[14'h28a0] = 8'hca;
s_mem_contents[14'h28a1] = 8'h10;
s_mem_contents[14'h28a2] = 8'he0;
s_mem_contents[14'h28a3] = 8'ha2;
s_mem_contents[14'h28a4] = 8'h03;
s_mem_contents[14'h28a5] = 8'ha9;
s_mem_contents[14'h28a6] = 8'h00;
s_mem_contents[14'h28a7] = 8'h48;
s_mem_contents[14'h28a8] = 8'hb5;
s_mem_contents[14'h28a9] = 8'h09;
s_mem_contents[14'h28aa] = 8'h9d;
s_mem_contents[14'h28ab] = 8'h03;
s_mem_contents[14'h28ac] = 8'h02;
s_mem_contents[14'h28ad] = 8'h28;
s_mem_contents[14'h28ae] = 8'h5e;
s_mem_contents[14'h28af] = 8'h03;
s_mem_contents[14'h28b0] = 8'h02;
s_mem_contents[14'h28b1] = 8'h08;
s_mem_contents[14'h28b2] = 8'hbd;
s_mem_contents[14'h28b3] = 8'h03;
s_mem_contents[14'h28b4] = 8'h02;
s_mem_contents[14'h28b5] = 8'hdd;
s_mem_contents[14'h28b6] = 8'h28;
s_mem_contents[14'h28b7] = 8'h02;
s_mem_contents[14'h28b8] = 8'hd0;
s_mem_contents[14'h28b9] = 8'hfe;
s_mem_contents[14'h28ba] = 8'h68;
s_mem_contents[14'h28bb] = 8'h49;
s_mem_contents[14'h28bc] = 8'h30;
s_mem_contents[14'h28bd] = 8'hdd;
s_mem_contents[14'h28be] = 8'h38;
s_mem_contents[14'h28bf] = 8'h02;
s_mem_contents[14'h28c0] = 8'hd0;
s_mem_contents[14'h28c1] = 8'hfe;
s_mem_contents[14'h28c2] = 8'hca;
s_mem_contents[14'h28c3] = 8'h10;
s_mem_contents[14'h28c4] = 8'he0;
s_mem_contents[14'h28c5] = 8'ha2;
s_mem_contents[14'h28c6] = 8'h03;
s_mem_contents[14'h28c7] = 8'ha9;
s_mem_contents[14'h28c8] = 8'hff;
s_mem_contents[14'h28c9] = 8'h48;
s_mem_contents[14'h28ca] = 8'hb5;
s_mem_contents[14'h28cb] = 8'h09;
s_mem_contents[14'h28cc] = 8'h9d;
s_mem_contents[14'h28cd] = 8'h03;
s_mem_contents[14'h28ce] = 8'h02;
s_mem_contents[14'h28cf] = 8'h28;
s_mem_contents[14'h28d0] = 8'h5e;
s_mem_contents[14'h28d1] = 8'h03;
s_mem_contents[14'h28d2] = 8'h02;
s_mem_contents[14'h28d3] = 8'h08;
s_mem_contents[14'h28d4] = 8'hbd;
s_mem_contents[14'h28d5] = 8'h03;
s_mem_contents[14'h28d6] = 8'h02;
s_mem_contents[14'h28d7] = 8'hdd;
s_mem_contents[14'h28d8] = 8'h28;
s_mem_contents[14'h28d9] = 8'h02;
s_mem_contents[14'h28da] = 8'hd0;
s_mem_contents[14'h28db] = 8'hfe;
s_mem_contents[14'h28dc] = 8'h68;
s_mem_contents[14'h28dd] = 8'h49;
s_mem_contents[14'h28de] = 8'h7c;
s_mem_contents[14'h28df] = 8'hdd;
s_mem_contents[14'h28e0] = 8'h38;
s_mem_contents[14'h28e1] = 8'h02;
s_mem_contents[14'h28e2] = 8'hd0;
s_mem_contents[14'h28e3] = 8'hfe;
s_mem_contents[14'h28e4] = 8'hca;
s_mem_contents[14'h28e5] = 8'h10;
s_mem_contents[14'h28e6] = 8'he0;
s_mem_contents[14'h28e7] = 8'ha2;
s_mem_contents[14'h28e8] = 8'h03;
s_mem_contents[14'h28e9] = 8'ha9;
s_mem_contents[14'h28ea] = 8'h00;
s_mem_contents[14'h28eb] = 8'h48;
s_mem_contents[14'h28ec] = 8'hb5;
s_mem_contents[14'h28ed] = 8'h09;
s_mem_contents[14'h28ee] = 8'h9d;
s_mem_contents[14'h28ef] = 8'h03;
s_mem_contents[14'h28f0] = 8'h02;
s_mem_contents[14'h28f1] = 8'h28;
s_mem_contents[14'h28f2] = 8'h3e;
s_mem_contents[14'h28f3] = 8'h03;
s_mem_contents[14'h28f4] = 8'h02;
s_mem_contents[14'h28f5] = 8'h08;
s_mem_contents[14'h28f6] = 8'hbd;
s_mem_contents[14'h28f7] = 8'h03;
s_mem_contents[14'h28f8] = 8'h02;
s_mem_contents[14'h28f9] = 8'hdd;
s_mem_contents[14'h28fa] = 8'h20;
s_mem_contents[14'h28fb] = 8'h02;
s_mem_contents[14'h28fc] = 8'hd0;
s_mem_contents[14'h28fd] = 8'hfe;
s_mem_contents[14'h28fe] = 8'h68;
s_mem_contents[14'h28ff] = 8'h49;
s_mem_contents[14'h2900] = 8'h30;
s_mem_contents[14'h2901] = 8'hdd;
s_mem_contents[14'h2902] = 8'h30;
s_mem_contents[14'h2903] = 8'h02;
s_mem_contents[14'h2904] = 8'hd0;
s_mem_contents[14'h2905] = 8'hfe;
s_mem_contents[14'h2906] = 8'hca;
s_mem_contents[14'h2907] = 8'h10;
s_mem_contents[14'h2908] = 8'he0;
s_mem_contents[14'h2909] = 8'ha2;
s_mem_contents[14'h290a] = 8'h03;
s_mem_contents[14'h290b] = 8'ha9;
s_mem_contents[14'h290c] = 8'hfe;
s_mem_contents[14'h290d] = 8'h48;
s_mem_contents[14'h290e] = 8'hb5;
s_mem_contents[14'h290f] = 8'h09;
s_mem_contents[14'h2910] = 8'h9d;
s_mem_contents[14'h2911] = 8'h03;
s_mem_contents[14'h2912] = 8'h02;
s_mem_contents[14'h2913] = 8'h28;
s_mem_contents[14'h2914] = 8'h3e;
s_mem_contents[14'h2915] = 8'h03;
s_mem_contents[14'h2916] = 8'h02;
s_mem_contents[14'h2917] = 8'h08;
s_mem_contents[14'h2918] = 8'hbd;
s_mem_contents[14'h2919] = 8'h03;
s_mem_contents[14'h291a] = 8'h02;
s_mem_contents[14'h291b] = 8'hdd;
s_mem_contents[14'h291c] = 8'h20;
s_mem_contents[14'h291d] = 8'h02;
s_mem_contents[14'h291e] = 8'hd0;
s_mem_contents[14'h291f] = 8'hfe;
s_mem_contents[14'h2920] = 8'h68;
s_mem_contents[14'h2921] = 8'h49;
s_mem_contents[14'h2922] = 8'h7c;
s_mem_contents[14'h2923] = 8'hdd;
s_mem_contents[14'h2924] = 8'h30;
s_mem_contents[14'h2925] = 8'h02;
s_mem_contents[14'h2926] = 8'hd0;
s_mem_contents[14'h2927] = 8'hfe;
s_mem_contents[14'h2928] = 8'hca;
s_mem_contents[14'h2929] = 8'h10;
s_mem_contents[14'h292a] = 8'he0;
s_mem_contents[14'h292b] = 8'ha2;
s_mem_contents[14'h292c] = 8'h03;
s_mem_contents[14'h292d] = 8'ha9;
s_mem_contents[14'h292e] = 8'h01;
s_mem_contents[14'h292f] = 8'h48;
s_mem_contents[14'h2930] = 8'hb5;
s_mem_contents[14'h2931] = 8'h09;
s_mem_contents[14'h2932] = 8'h9d;
s_mem_contents[14'h2933] = 8'h03;
s_mem_contents[14'h2934] = 8'h02;
s_mem_contents[14'h2935] = 8'h28;
s_mem_contents[14'h2936] = 8'h3e;
s_mem_contents[14'h2937] = 8'h03;
s_mem_contents[14'h2938] = 8'h02;
s_mem_contents[14'h2939] = 8'h08;
s_mem_contents[14'h293a] = 8'hbd;
s_mem_contents[14'h293b] = 8'h03;
s_mem_contents[14'h293c] = 8'h02;
s_mem_contents[14'h293d] = 8'hdd;
s_mem_contents[14'h293e] = 8'h24;
s_mem_contents[14'h293f] = 8'h02;
s_mem_contents[14'h2940] = 8'hd0;
s_mem_contents[14'h2941] = 8'hfe;
s_mem_contents[14'h2942] = 8'h68;
s_mem_contents[14'h2943] = 8'h49;
s_mem_contents[14'h2944] = 8'h30;
s_mem_contents[14'h2945] = 8'hdd;
s_mem_contents[14'h2946] = 8'h34;
s_mem_contents[14'h2947] = 8'h02;
s_mem_contents[14'h2948] = 8'hd0;
s_mem_contents[14'h2949] = 8'hfe;
s_mem_contents[14'h294a] = 8'hca;
s_mem_contents[14'h294b] = 8'h10;
s_mem_contents[14'h294c] = 8'he0;
s_mem_contents[14'h294d] = 8'ha2;
s_mem_contents[14'h294e] = 8'h03;
s_mem_contents[14'h294f] = 8'ha9;
s_mem_contents[14'h2950] = 8'hff;
s_mem_contents[14'h2951] = 8'h48;
s_mem_contents[14'h2952] = 8'hb5;
s_mem_contents[14'h2953] = 8'h09;
s_mem_contents[14'h2954] = 8'h9d;
s_mem_contents[14'h2955] = 8'h03;
s_mem_contents[14'h2956] = 8'h02;
s_mem_contents[14'h2957] = 8'h28;
s_mem_contents[14'h2958] = 8'h3e;
s_mem_contents[14'h2959] = 8'h03;
s_mem_contents[14'h295a] = 8'h02;
s_mem_contents[14'h295b] = 8'h08;
s_mem_contents[14'h295c] = 8'hbd;
s_mem_contents[14'h295d] = 8'h03;
s_mem_contents[14'h295e] = 8'h02;
s_mem_contents[14'h295f] = 8'hdd;
s_mem_contents[14'h2960] = 8'h24;
s_mem_contents[14'h2961] = 8'h02;
s_mem_contents[14'h2962] = 8'hd0;
s_mem_contents[14'h2963] = 8'hfe;
s_mem_contents[14'h2964] = 8'h68;
s_mem_contents[14'h2965] = 8'h49;
s_mem_contents[14'h2966] = 8'h7c;
s_mem_contents[14'h2967] = 8'hdd;
s_mem_contents[14'h2968] = 8'h34;
s_mem_contents[14'h2969] = 8'h02;
s_mem_contents[14'h296a] = 8'hd0;
s_mem_contents[14'h296b] = 8'hfe;
s_mem_contents[14'h296c] = 8'hca;
s_mem_contents[14'h296d] = 8'h10;
s_mem_contents[14'h296e] = 8'he0;
s_mem_contents[14'h296f] = 8'ha2;
s_mem_contents[14'h2970] = 8'h03;
s_mem_contents[14'h2971] = 8'ha9;
s_mem_contents[14'h2972] = 8'h00;
s_mem_contents[14'h2973] = 8'h48;
s_mem_contents[14'h2974] = 8'hb5;
s_mem_contents[14'h2975] = 8'h09;
s_mem_contents[14'h2976] = 8'h9d;
s_mem_contents[14'h2977] = 8'h03;
s_mem_contents[14'h2978] = 8'h02;
s_mem_contents[14'h2979] = 8'h28;
s_mem_contents[14'h297a] = 8'h7e;
s_mem_contents[14'h297b] = 8'h03;
s_mem_contents[14'h297c] = 8'h02;
s_mem_contents[14'h297d] = 8'h08;
s_mem_contents[14'h297e] = 8'hbd;
s_mem_contents[14'h297f] = 8'h03;
s_mem_contents[14'h2980] = 8'h02;
s_mem_contents[14'h2981] = 8'hdd;
s_mem_contents[14'h2982] = 8'h28;
s_mem_contents[14'h2983] = 8'h02;
s_mem_contents[14'h2984] = 8'hd0;
s_mem_contents[14'h2985] = 8'hfe;
s_mem_contents[14'h2986] = 8'h68;
s_mem_contents[14'h2987] = 8'h49;
s_mem_contents[14'h2988] = 8'h30;
s_mem_contents[14'h2989] = 8'hdd;
s_mem_contents[14'h298a] = 8'h38;
s_mem_contents[14'h298b] = 8'h02;
s_mem_contents[14'h298c] = 8'hd0;
s_mem_contents[14'h298d] = 8'hfe;
s_mem_contents[14'h298e] = 8'hca;
s_mem_contents[14'h298f] = 8'h10;
s_mem_contents[14'h2990] = 8'he0;
s_mem_contents[14'h2991] = 8'ha2;
s_mem_contents[14'h2992] = 8'h03;
s_mem_contents[14'h2993] = 8'ha9;
s_mem_contents[14'h2994] = 8'hfe;
s_mem_contents[14'h2995] = 8'h48;
s_mem_contents[14'h2996] = 8'hb5;
s_mem_contents[14'h2997] = 8'h09;
s_mem_contents[14'h2998] = 8'h9d;
s_mem_contents[14'h2999] = 8'h03;
s_mem_contents[14'h299a] = 8'h02;
s_mem_contents[14'h299b] = 8'h28;
s_mem_contents[14'h299c] = 8'h7e;
s_mem_contents[14'h299d] = 8'h03;
s_mem_contents[14'h299e] = 8'h02;
s_mem_contents[14'h299f] = 8'h08;
s_mem_contents[14'h29a0] = 8'hbd;
s_mem_contents[14'h29a1] = 8'h03;
s_mem_contents[14'h29a2] = 8'h02;
s_mem_contents[14'h29a3] = 8'hdd;
s_mem_contents[14'h29a4] = 8'h28;
s_mem_contents[14'h29a5] = 8'h02;
s_mem_contents[14'h29a6] = 8'hd0;
s_mem_contents[14'h29a7] = 8'hfe;
s_mem_contents[14'h29a8] = 8'h68;
s_mem_contents[14'h29a9] = 8'h49;
s_mem_contents[14'h29aa] = 8'h7c;
s_mem_contents[14'h29ab] = 8'hdd;
s_mem_contents[14'h29ac] = 8'h38;
s_mem_contents[14'h29ad] = 8'h02;
s_mem_contents[14'h29ae] = 8'hd0;
s_mem_contents[14'h29af] = 8'hfe;
s_mem_contents[14'h29b0] = 8'hca;
s_mem_contents[14'h29b1] = 8'h10;
s_mem_contents[14'h29b2] = 8'he0;
s_mem_contents[14'h29b3] = 8'ha2;
s_mem_contents[14'h29b4] = 8'h03;
s_mem_contents[14'h29b5] = 8'ha9;
s_mem_contents[14'h29b6] = 8'h01;
s_mem_contents[14'h29b7] = 8'h48;
s_mem_contents[14'h29b8] = 8'hb5;
s_mem_contents[14'h29b9] = 8'h09;
s_mem_contents[14'h29ba] = 8'h9d;
s_mem_contents[14'h29bb] = 8'h03;
s_mem_contents[14'h29bc] = 8'h02;
s_mem_contents[14'h29bd] = 8'h28;
s_mem_contents[14'h29be] = 8'h7e;
s_mem_contents[14'h29bf] = 8'h03;
s_mem_contents[14'h29c0] = 8'h02;
s_mem_contents[14'h29c1] = 8'h08;
s_mem_contents[14'h29c2] = 8'hbd;
s_mem_contents[14'h29c3] = 8'h03;
s_mem_contents[14'h29c4] = 8'h02;
s_mem_contents[14'h29c5] = 8'hdd;
s_mem_contents[14'h29c6] = 8'h2c;
s_mem_contents[14'h29c7] = 8'h02;
s_mem_contents[14'h29c8] = 8'hd0;
s_mem_contents[14'h29c9] = 8'hfe;
s_mem_contents[14'h29ca] = 8'h68;
s_mem_contents[14'h29cb] = 8'h49;
s_mem_contents[14'h29cc] = 8'h30;
s_mem_contents[14'h29cd] = 8'hdd;
s_mem_contents[14'h29ce] = 8'h3c;
s_mem_contents[14'h29cf] = 8'h02;
s_mem_contents[14'h29d0] = 8'hd0;
s_mem_contents[14'h29d1] = 8'hfe;
s_mem_contents[14'h29d2] = 8'hca;
s_mem_contents[14'h29d3] = 8'h10;
s_mem_contents[14'h29d4] = 8'he0;
s_mem_contents[14'h29d5] = 8'ha2;
s_mem_contents[14'h29d6] = 8'h03;
s_mem_contents[14'h29d7] = 8'ha9;
s_mem_contents[14'h29d8] = 8'hff;
s_mem_contents[14'h29d9] = 8'h48;
s_mem_contents[14'h29da] = 8'hb5;
s_mem_contents[14'h29db] = 8'h09;
s_mem_contents[14'h29dc] = 8'h9d;
s_mem_contents[14'h29dd] = 8'h03;
s_mem_contents[14'h29de] = 8'h02;
s_mem_contents[14'h29df] = 8'h28;
s_mem_contents[14'h29e0] = 8'h7e;
s_mem_contents[14'h29e1] = 8'h03;
s_mem_contents[14'h29e2] = 8'h02;
s_mem_contents[14'h29e3] = 8'h08;
s_mem_contents[14'h29e4] = 8'hbd;
s_mem_contents[14'h29e5] = 8'h03;
s_mem_contents[14'h29e6] = 8'h02;
s_mem_contents[14'h29e7] = 8'hdd;
s_mem_contents[14'h29e8] = 8'h2c;
s_mem_contents[14'h29e9] = 8'h02;
s_mem_contents[14'h29ea] = 8'hd0;
s_mem_contents[14'h29eb] = 8'hfe;
s_mem_contents[14'h29ec] = 8'h68;
s_mem_contents[14'h29ed] = 8'h49;
s_mem_contents[14'h29ee] = 8'h7c;
s_mem_contents[14'h29ef] = 8'hdd;
s_mem_contents[14'h29f0] = 8'h3c;
s_mem_contents[14'h29f1] = 8'h02;
s_mem_contents[14'h29f2] = 8'hd0;
s_mem_contents[14'h29f3] = 8'hfe;
s_mem_contents[14'h29f4] = 8'hca;
s_mem_contents[14'h29f5] = 8'h10;
s_mem_contents[14'h29f6] = 8'he0;
s_mem_contents[14'h29f7] = 8'had;
s_mem_contents[14'h29f8] = 8'h00;
s_mem_contents[14'h29f9] = 8'h02;
s_mem_contents[14'h29fa] = 8'hc9;
s_mem_contents[14'h29fb] = 8'h21;
s_mem_contents[14'h29fc] = 8'hd0;
s_mem_contents[14'h29fd] = 8'hfe;
s_mem_contents[14'h29fe] = 8'ha9;
s_mem_contents[14'h29ff] = 8'h22;
s_mem_contents[14'h2a00] = 8'h8d;
s_mem_contents[14'h2a01] = 8'h00;
s_mem_contents[14'h2a02] = 8'h02;
s_mem_contents[14'h2a03] = 8'ha2;
s_mem_contents[14'h2a04] = 8'h00;
s_mem_contents[14'h2a05] = 8'ha9;
s_mem_contents[14'h2a06] = 8'h7e;
s_mem_contents[14'h2a07] = 8'h85;
s_mem_contents[14'h2a08] = 8'h02;
s_mem_contents[14'h2a09] = 8'ha9;
s_mem_contents[14'h2a0a] = 8'h00;
s_mem_contents[14'h2a0b] = 8'h48;
s_mem_contents[14'h2a0c] = 8'h28;
s_mem_contents[14'h2a0d] = 8'he6;
s_mem_contents[14'h2a0e] = 8'h02;
s_mem_contents[14'h2a0f] = 8'h08;
s_mem_contents[14'h2a10] = 8'ha5;
s_mem_contents[14'h2a11] = 8'h02;
s_mem_contents[14'h2a12] = 8'hdd;
s_mem_contents[14'h2a13] = 8'h40;
s_mem_contents[14'h2a14] = 8'h02;
s_mem_contents[14'h2a15] = 8'hd0;
s_mem_contents[14'h2a16] = 8'hfe;
s_mem_contents[14'h2a17] = 8'h68;
s_mem_contents[14'h2a18] = 8'h49;
s_mem_contents[14'h2a19] = 8'h30;
s_mem_contents[14'h2a1a] = 8'hdd;
s_mem_contents[14'h2a1b] = 8'h45;
s_mem_contents[14'h2a1c] = 8'h02;
s_mem_contents[14'h2a1d] = 8'hd0;
s_mem_contents[14'h2a1e] = 8'hfe;
s_mem_contents[14'h2a1f] = 8'he8;
s_mem_contents[14'h2a20] = 8'he0;
s_mem_contents[14'h2a21] = 8'h02;
s_mem_contents[14'h2a22] = 8'hd0;
s_mem_contents[14'h2a23] = 8'h04;
s_mem_contents[14'h2a24] = 8'ha9;
s_mem_contents[14'h2a25] = 8'hfe;
s_mem_contents[14'h2a26] = 8'h85;
s_mem_contents[14'h2a27] = 8'h02;
s_mem_contents[14'h2a28] = 8'he0;
s_mem_contents[14'h2a29] = 8'h05;
s_mem_contents[14'h2a2a] = 8'hd0;
s_mem_contents[14'h2a2b] = 8'hdd;
s_mem_contents[14'h2a2c] = 8'hca;
s_mem_contents[14'h2a2d] = 8'he6;
s_mem_contents[14'h2a2e] = 8'h02;
s_mem_contents[14'h2a2f] = 8'ha9;
s_mem_contents[14'h2a30] = 8'h00;
s_mem_contents[14'h2a31] = 8'h48;
s_mem_contents[14'h2a32] = 8'h28;
s_mem_contents[14'h2a33] = 8'hc6;
s_mem_contents[14'h2a34] = 8'h02;
s_mem_contents[14'h2a35] = 8'h08;
s_mem_contents[14'h2a36] = 8'ha5;
s_mem_contents[14'h2a37] = 8'h02;
s_mem_contents[14'h2a38] = 8'hdd;
s_mem_contents[14'h2a39] = 8'h40;
s_mem_contents[14'h2a3a] = 8'h02;
s_mem_contents[14'h2a3b] = 8'hd0;
s_mem_contents[14'h2a3c] = 8'hfe;
s_mem_contents[14'h2a3d] = 8'h68;
s_mem_contents[14'h2a3e] = 8'h49;
s_mem_contents[14'h2a3f] = 8'h30;
s_mem_contents[14'h2a40] = 8'hdd;
s_mem_contents[14'h2a41] = 8'h45;
s_mem_contents[14'h2a42] = 8'h02;
s_mem_contents[14'h2a43] = 8'hd0;
s_mem_contents[14'h2a44] = 8'hfe;
s_mem_contents[14'h2a45] = 8'hca;
s_mem_contents[14'h2a46] = 8'h30;
s_mem_contents[14'h2a47] = 8'h0a;
s_mem_contents[14'h2a48] = 8'he0;
s_mem_contents[14'h2a49] = 8'h01;
s_mem_contents[14'h2a4a] = 8'hd0;
s_mem_contents[14'h2a4b] = 8'he3;
s_mem_contents[14'h2a4c] = 8'ha9;
s_mem_contents[14'h2a4d] = 8'h81;
s_mem_contents[14'h2a4e] = 8'h85;
s_mem_contents[14'h2a4f] = 8'h02;
s_mem_contents[14'h2a50] = 8'hd0;
s_mem_contents[14'h2a51] = 8'hdd;
s_mem_contents[14'h2a52] = 8'ha2;
s_mem_contents[14'h2a53] = 8'h00;
s_mem_contents[14'h2a54] = 8'ha9;
s_mem_contents[14'h2a55] = 8'h7e;
s_mem_contents[14'h2a56] = 8'h85;
s_mem_contents[14'h2a57] = 8'h02;
s_mem_contents[14'h2a58] = 8'ha9;
s_mem_contents[14'h2a59] = 8'hff;
s_mem_contents[14'h2a5a] = 8'h48;
s_mem_contents[14'h2a5b] = 8'h28;
s_mem_contents[14'h2a5c] = 8'he6;
s_mem_contents[14'h2a5d] = 8'h02;
s_mem_contents[14'h2a5e] = 8'h08;
s_mem_contents[14'h2a5f] = 8'ha5;
s_mem_contents[14'h2a60] = 8'h02;
s_mem_contents[14'h2a61] = 8'hdd;
s_mem_contents[14'h2a62] = 8'h40;
s_mem_contents[14'h2a63] = 8'h02;
s_mem_contents[14'h2a64] = 8'hd0;
s_mem_contents[14'h2a65] = 8'hfe;
s_mem_contents[14'h2a66] = 8'h68;
s_mem_contents[14'h2a67] = 8'h49;
s_mem_contents[14'h2a68] = 8'h7d;
s_mem_contents[14'h2a69] = 8'hdd;
s_mem_contents[14'h2a6a] = 8'h45;
s_mem_contents[14'h2a6b] = 8'h02;
s_mem_contents[14'h2a6c] = 8'hd0;
s_mem_contents[14'h2a6d] = 8'hfe;
s_mem_contents[14'h2a6e] = 8'he8;
s_mem_contents[14'h2a6f] = 8'he0;
s_mem_contents[14'h2a70] = 8'h02;
s_mem_contents[14'h2a71] = 8'hd0;
s_mem_contents[14'h2a72] = 8'h04;
s_mem_contents[14'h2a73] = 8'ha9;
s_mem_contents[14'h2a74] = 8'hfe;
s_mem_contents[14'h2a75] = 8'h85;
s_mem_contents[14'h2a76] = 8'h02;
s_mem_contents[14'h2a77] = 8'he0;
s_mem_contents[14'h2a78] = 8'h05;
s_mem_contents[14'h2a79] = 8'hd0;
s_mem_contents[14'h2a7a] = 8'hdd;
s_mem_contents[14'h2a7b] = 8'hca;
s_mem_contents[14'h2a7c] = 8'he6;
s_mem_contents[14'h2a7d] = 8'h02;
s_mem_contents[14'h2a7e] = 8'ha9;
s_mem_contents[14'h2a7f] = 8'hff;
s_mem_contents[14'h2a80] = 8'h48;
s_mem_contents[14'h2a81] = 8'h28;
s_mem_contents[14'h2a82] = 8'hc6;
s_mem_contents[14'h2a83] = 8'h02;
s_mem_contents[14'h2a84] = 8'h08;
s_mem_contents[14'h2a85] = 8'ha5;
s_mem_contents[14'h2a86] = 8'h02;
s_mem_contents[14'h2a87] = 8'hdd;
s_mem_contents[14'h2a88] = 8'h40;
s_mem_contents[14'h2a89] = 8'h02;
s_mem_contents[14'h2a8a] = 8'hd0;
s_mem_contents[14'h2a8b] = 8'hfe;
s_mem_contents[14'h2a8c] = 8'h68;
s_mem_contents[14'h2a8d] = 8'h49;
s_mem_contents[14'h2a8e] = 8'h7d;
s_mem_contents[14'h2a8f] = 8'hdd;
s_mem_contents[14'h2a90] = 8'h45;
s_mem_contents[14'h2a91] = 8'h02;
s_mem_contents[14'h2a92] = 8'hd0;
s_mem_contents[14'h2a93] = 8'hfe;
s_mem_contents[14'h2a94] = 8'hca;
s_mem_contents[14'h2a95] = 8'h30;
s_mem_contents[14'h2a96] = 8'h0a;
s_mem_contents[14'h2a97] = 8'he0;
s_mem_contents[14'h2a98] = 8'h01;
s_mem_contents[14'h2a99] = 8'hd0;
s_mem_contents[14'h2a9a] = 8'he3;
s_mem_contents[14'h2a9b] = 8'ha9;
s_mem_contents[14'h2a9c] = 8'h81;
s_mem_contents[14'h2a9d] = 8'h85;
s_mem_contents[14'h2a9e] = 8'h02;
s_mem_contents[14'h2a9f] = 8'hd0;
s_mem_contents[14'h2aa0] = 8'hdd;
s_mem_contents[14'h2aa1] = 8'had;
s_mem_contents[14'h2aa2] = 8'h00;
s_mem_contents[14'h2aa3] = 8'h02;
s_mem_contents[14'h2aa4] = 8'hc9;
s_mem_contents[14'h2aa5] = 8'h22;
s_mem_contents[14'h2aa6] = 8'hd0;
s_mem_contents[14'h2aa7] = 8'hfe;
s_mem_contents[14'h2aa8] = 8'ha9;
s_mem_contents[14'h2aa9] = 8'h23;
s_mem_contents[14'h2aaa] = 8'h8d;
s_mem_contents[14'h2aab] = 8'h00;
s_mem_contents[14'h2aac] = 8'h02;
s_mem_contents[14'h2aad] = 8'ha2;
s_mem_contents[14'h2aae] = 8'h00;
s_mem_contents[14'h2aaf] = 8'ha9;
s_mem_contents[14'h2ab0] = 8'h7e;
s_mem_contents[14'h2ab1] = 8'h8d;
s_mem_contents[14'h2ab2] = 8'h03;
s_mem_contents[14'h2ab3] = 8'h02;
s_mem_contents[14'h2ab4] = 8'ha9;
s_mem_contents[14'h2ab5] = 8'h00;
s_mem_contents[14'h2ab6] = 8'h48;
s_mem_contents[14'h2ab7] = 8'h28;
s_mem_contents[14'h2ab8] = 8'hee;
s_mem_contents[14'h2ab9] = 8'h03;
s_mem_contents[14'h2aba] = 8'h02;
s_mem_contents[14'h2abb] = 8'h08;
s_mem_contents[14'h2abc] = 8'had;
s_mem_contents[14'h2abd] = 8'h03;
s_mem_contents[14'h2abe] = 8'h02;
s_mem_contents[14'h2abf] = 8'hdd;
s_mem_contents[14'h2ac0] = 8'h40;
s_mem_contents[14'h2ac1] = 8'h02;
s_mem_contents[14'h2ac2] = 8'hd0;
s_mem_contents[14'h2ac3] = 8'hfe;
s_mem_contents[14'h2ac4] = 8'h68;
s_mem_contents[14'h2ac5] = 8'h49;
s_mem_contents[14'h2ac6] = 8'h30;
s_mem_contents[14'h2ac7] = 8'hdd;
s_mem_contents[14'h2ac8] = 8'h45;
s_mem_contents[14'h2ac9] = 8'h02;
s_mem_contents[14'h2aca] = 8'hd0;
s_mem_contents[14'h2acb] = 8'hfe;
s_mem_contents[14'h2acc] = 8'he8;
s_mem_contents[14'h2acd] = 8'he0;
s_mem_contents[14'h2ace] = 8'h02;
s_mem_contents[14'h2acf] = 8'hd0;
s_mem_contents[14'h2ad0] = 8'h05;
s_mem_contents[14'h2ad1] = 8'ha9;
s_mem_contents[14'h2ad2] = 8'hfe;
s_mem_contents[14'h2ad3] = 8'h8d;
s_mem_contents[14'h2ad4] = 8'h03;
s_mem_contents[14'h2ad5] = 8'h02;
s_mem_contents[14'h2ad6] = 8'he0;
s_mem_contents[14'h2ad7] = 8'h05;
s_mem_contents[14'h2ad8] = 8'hd0;
s_mem_contents[14'h2ad9] = 8'hda;
s_mem_contents[14'h2ada] = 8'hca;
s_mem_contents[14'h2adb] = 8'hee;
s_mem_contents[14'h2adc] = 8'h03;
s_mem_contents[14'h2add] = 8'h02;
s_mem_contents[14'h2ade] = 8'ha9;
s_mem_contents[14'h2adf] = 8'h00;
s_mem_contents[14'h2ae0] = 8'h48;
s_mem_contents[14'h2ae1] = 8'h28;
s_mem_contents[14'h2ae2] = 8'hce;
s_mem_contents[14'h2ae3] = 8'h03;
s_mem_contents[14'h2ae4] = 8'h02;
s_mem_contents[14'h2ae5] = 8'h08;
s_mem_contents[14'h2ae6] = 8'had;
s_mem_contents[14'h2ae7] = 8'h03;
s_mem_contents[14'h2ae8] = 8'h02;
s_mem_contents[14'h2ae9] = 8'hdd;
s_mem_contents[14'h2aea] = 8'h40;
s_mem_contents[14'h2aeb] = 8'h02;
s_mem_contents[14'h2aec] = 8'hd0;
s_mem_contents[14'h2aed] = 8'hfe;
s_mem_contents[14'h2aee] = 8'h68;
s_mem_contents[14'h2aef] = 8'h49;
s_mem_contents[14'h2af0] = 8'h30;
s_mem_contents[14'h2af1] = 8'hdd;
s_mem_contents[14'h2af2] = 8'h45;
s_mem_contents[14'h2af3] = 8'h02;
s_mem_contents[14'h2af4] = 8'hd0;
s_mem_contents[14'h2af5] = 8'hfe;
s_mem_contents[14'h2af6] = 8'hca;
s_mem_contents[14'h2af7] = 8'h30;
s_mem_contents[14'h2af8] = 8'h0b;
s_mem_contents[14'h2af9] = 8'he0;
s_mem_contents[14'h2afa] = 8'h01;
s_mem_contents[14'h2afb] = 8'hd0;
s_mem_contents[14'h2afc] = 8'he1;
s_mem_contents[14'h2afd] = 8'ha9;
s_mem_contents[14'h2afe] = 8'h81;
s_mem_contents[14'h2aff] = 8'h8d;
s_mem_contents[14'h2b00] = 8'h03;
s_mem_contents[14'h2b01] = 8'h02;
s_mem_contents[14'h2b02] = 8'hd0;
s_mem_contents[14'h2b03] = 8'hda;
s_mem_contents[14'h2b04] = 8'ha2;
s_mem_contents[14'h2b05] = 8'h00;
s_mem_contents[14'h2b06] = 8'ha9;
s_mem_contents[14'h2b07] = 8'h7e;
s_mem_contents[14'h2b08] = 8'h8d;
s_mem_contents[14'h2b09] = 8'h03;
s_mem_contents[14'h2b0a] = 8'h02;
s_mem_contents[14'h2b0b] = 8'ha9;
s_mem_contents[14'h2b0c] = 8'hff;
s_mem_contents[14'h2b0d] = 8'h48;
s_mem_contents[14'h2b0e] = 8'h28;
s_mem_contents[14'h2b0f] = 8'hee;
s_mem_contents[14'h2b10] = 8'h03;
s_mem_contents[14'h2b11] = 8'h02;
s_mem_contents[14'h2b12] = 8'h08;
s_mem_contents[14'h2b13] = 8'had;
s_mem_contents[14'h2b14] = 8'h03;
s_mem_contents[14'h2b15] = 8'h02;
s_mem_contents[14'h2b16] = 8'hdd;
s_mem_contents[14'h2b17] = 8'h40;
s_mem_contents[14'h2b18] = 8'h02;
s_mem_contents[14'h2b19] = 8'hd0;
s_mem_contents[14'h2b1a] = 8'hfe;
s_mem_contents[14'h2b1b] = 8'h68;
s_mem_contents[14'h2b1c] = 8'h49;
s_mem_contents[14'h2b1d] = 8'h7d;
s_mem_contents[14'h2b1e] = 8'hdd;
s_mem_contents[14'h2b1f] = 8'h45;
s_mem_contents[14'h2b20] = 8'h02;
s_mem_contents[14'h2b21] = 8'hd0;
s_mem_contents[14'h2b22] = 8'hfe;
s_mem_contents[14'h2b23] = 8'he8;
s_mem_contents[14'h2b24] = 8'he0;
s_mem_contents[14'h2b25] = 8'h02;
s_mem_contents[14'h2b26] = 8'hd0;
s_mem_contents[14'h2b27] = 8'h05;
s_mem_contents[14'h2b28] = 8'ha9;
s_mem_contents[14'h2b29] = 8'hfe;
s_mem_contents[14'h2b2a] = 8'h8d;
s_mem_contents[14'h2b2b] = 8'h03;
s_mem_contents[14'h2b2c] = 8'h02;
s_mem_contents[14'h2b2d] = 8'he0;
s_mem_contents[14'h2b2e] = 8'h05;
s_mem_contents[14'h2b2f] = 8'hd0;
s_mem_contents[14'h2b30] = 8'hda;
s_mem_contents[14'h2b31] = 8'hca;
s_mem_contents[14'h2b32] = 8'hee;
s_mem_contents[14'h2b33] = 8'h03;
s_mem_contents[14'h2b34] = 8'h02;
s_mem_contents[14'h2b35] = 8'ha9;
s_mem_contents[14'h2b36] = 8'hff;
s_mem_contents[14'h2b37] = 8'h48;
s_mem_contents[14'h2b38] = 8'h28;
s_mem_contents[14'h2b39] = 8'hce;
s_mem_contents[14'h2b3a] = 8'h03;
s_mem_contents[14'h2b3b] = 8'h02;
s_mem_contents[14'h2b3c] = 8'h08;
s_mem_contents[14'h2b3d] = 8'had;
s_mem_contents[14'h2b3e] = 8'h03;
s_mem_contents[14'h2b3f] = 8'h02;
s_mem_contents[14'h2b40] = 8'hdd;
s_mem_contents[14'h2b41] = 8'h40;
s_mem_contents[14'h2b42] = 8'h02;
s_mem_contents[14'h2b43] = 8'hd0;
s_mem_contents[14'h2b44] = 8'hfe;
s_mem_contents[14'h2b45] = 8'h68;
s_mem_contents[14'h2b46] = 8'h49;
s_mem_contents[14'h2b47] = 8'h7d;
s_mem_contents[14'h2b48] = 8'hdd;
s_mem_contents[14'h2b49] = 8'h45;
s_mem_contents[14'h2b4a] = 8'h02;
s_mem_contents[14'h2b4b] = 8'hd0;
s_mem_contents[14'h2b4c] = 8'hfe;
s_mem_contents[14'h2b4d] = 8'hca;
s_mem_contents[14'h2b4e] = 8'h30;
s_mem_contents[14'h2b4f] = 8'h0b;
s_mem_contents[14'h2b50] = 8'he0;
s_mem_contents[14'h2b51] = 8'h01;
s_mem_contents[14'h2b52] = 8'hd0;
s_mem_contents[14'h2b53] = 8'he1;
s_mem_contents[14'h2b54] = 8'ha9;
s_mem_contents[14'h2b55] = 8'h81;
s_mem_contents[14'h2b56] = 8'h8d;
s_mem_contents[14'h2b57] = 8'h03;
s_mem_contents[14'h2b58] = 8'h02;
s_mem_contents[14'h2b59] = 8'hd0;
s_mem_contents[14'h2b5a] = 8'hda;
s_mem_contents[14'h2b5b] = 8'had;
s_mem_contents[14'h2b5c] = 8'h00;
s_mem_contents[14'h2b5d] = 8'h02;
s_mem_contents[14'h2b5e] = 8'hc9;
s_mem_contents[14'h2b5f] = 8'h23;
s_mem_contents[14'h2b60] = 8'hd0;
s_mem_contents[14'h2b61] = 8'hfe;
s_mem_contents[14'h2b62] = 8'ha9;
s_mem_contents[14'h2b63] = 8'h24;
s_mem_contents[14'h2b64] = 8'h8d;
s_mem_contents[14'h2b65] = 8'h00;
s_mem_contents[14'h2b66] = 8'h02;
s_mem_contents[14'h2b67] = 8'ha2;
s_mem_contents[14'h2b68] = 8'h00;
s_mem_contents[14'h2b69] = 8'ha9;
s_mem_contents[14'h2b6a] = 8'h7e;
s_mem_contents[14'h2b6b] = 8'h95;
s_mem_contents[14'h2b6c] = 8'h02;
s_mem_contents[14'h2b6d] = 8'ha9;
s_mem_contents[14'h2b6e] = 8'h00;
s_mem_contents[14'h2b6f] = 8'h48;
s_mem_contents[14'h2b70] = 8'h28;
s_mem_contents[14'h2b71] = 8'hf6;
s_mem_contents[14'h2b72] = 8'h02;
s_mem_contents[14'h2b73] = 8'h08;
s_mem_contents[14'h2b74] = 8'hb5;
s_mem_contents[14'h2b75] = 8'h02;
s_mem_contents[14'h2b76] = 8'hdd;
s_mem_contents[14'h2b77] = 8'h40;
s_mem_contents[14'h2b78] = 8'h02;
s_mem_contents[14'h2b79] = 8'hd0;
s_mem_contents[14'h2b7a] = 8'hfe;
s_mem_contents[14'h2b7b] = 8'h68;
s_mem_contents[14'h2b7c] = 8'h49;
s_mem_contents[14'h2b7d] = 8'h30;
s_mem_contents[14'h2b7e] = 8'hdd;
s_mem_contents[14'h2b7f] = 8'h45;
s_mem_contents[14'h2b80] = 8'h02;
s_mem_contents[14'h2b81] = 8'hd0;
s_mem_contents[14'h2b82] = 8'hfe;
s_mem_contents[14'h2b83] = 8'hb5;
s_mem_contents[14'h2b84] = 8'h02;
s_mem_contents[14'h2b85] = 8'he8;
s_mem_contents[14'h2b86] = 8'he0;
s_mem_contents[14'h2b87] = 8'h02;
s_mem_contents[14'h2b88] = 8'hd0;
s_mem_contents[14'h2b89] = 8'h02;
s_mem_contents[14'h2b8a] = 8'ha9;
s_mem_contents[14'h2b8b] = 8'hfe;
s_mem_contents[14'h2b8c] = 8'he0;
s_mem_contents[14'h2b8d] = 8'h05;
s_mem_contents[14'h2b8e] = 8'hd0;
s_mem_contents[14'h2b8f] = 8'hdb;
s_mem_contents[14'h2b90] = 8'hca;
s_mem_contents[14'h2b91] = 8'ha9;
s_mem_contents[14'h2b92] = 8'h02;
s_mem_contents[14'h2b93] = 8'h95;
s_mem_contents[14'h2b94] = 8'h02;
s_mem_contents[14'h2b95] = 8'ha9;
s_mem_contents[14'h2b96] = 8'h00;
s_mem_contents[14'h2b97] = 8'h48;
s_mem_contents[14'h2b98] = 8'h28;
s_mem_contents[14'h2b99] = 8'hd6;
s_mem_contents[14'h2b9a] = 8'h02;
s_mem_contents[14'h2b9b] = 8'h08;
s_mem_contents[14'h2b9c] = 8'hb5;
s_mem_contents[14'h2b9d] = 8'h02;
s_mem_contents[14'h2b9e] = 8'hdd;
s_mem_contents[14'h2b9f] = 8'h40;
s_mem_contents[14'h2ba0] = 8'h02;
s_mem_contents[14'h2ba1] = 8'hd0;
s_mem_contents[14'h2ba2] = 8'hfe;
s_mem_contents[14'h2ba3] = 8'h68;
s_mem_contents[14'h2ba4] = 8'h49;
s_mem_contents[14'h2ba5] = 8'h30;
s_mem_contents[14'h2ba6] = 8'hdd;
s_mem_contents[14'h2ba7] = 8'h45;
s_mem_contents[14'h2ba8] = 8'h02;
s_mem_contents[14'h2ba9] = 8'hd0;
s_mem_contents[14'h2baa] = 8'hfe;
s_mem_contents[14'h2bab] = 8'hb5;
s_mem_contents[14'h2bac] = 8'h02;
s_mem_contents[14'h2bad] = 8'hca;
s_mem_contents[14'h2bae] = 8'h30;
s_mem_contents[14'h2baf] = 8'h08;
s_mem_contents[14'h2bb0] = 8'he0;
s_mem_contents[14'h2bb1] = 8'h01;
s_mem_contents[14'h2bb2] = 8'hd0;
s_mem_contents[14'h2bb3] = 8'hdf;
s_mem_contents[14'h2bb4] = 8'ha9;
s_mem_contents[14'h2bb5] = 8'h81;
s_mem_contents[14'h2bb6] = 8'hd0;
s_mem_contents[14'h2bb7] = 8'hdb;
s_mem_contents[14'h2bb8] = 8'ha2;
s_mem_contents[14'h2bb9] = 8'h00;
s_mem_contents[14'h2bba] = 8'ha9;
s_mem_contents[14'h2bbb] = 8'h7e;
s_mem_contents[14'h2bbc] = 8'h95;
s_mem_contents[14'h2bbd] = 8'h02;
s_mem_contents[14'h2bbe] = 8'ha9;
s_mem_contents[14'h2bbf] = 8'hff;
s_mem_contents[14'h2bc0] = 8'h48;
s_mem_contents[14'h2bc1] = 8'h28;
s_mem_contents[14'h2bc2] = 8'hf6;
s_mem_contents[14'h2bc3] = 8'h02;
s_mem_contents[14'h2bc4] = 8'h08;
s_mem_contents[14'h2bc5] = 8'hb5;
s_mem_contents[14'h2bc6] = 8'h02;
s_mem_contents[14'h2bc7] = 8'hdd;
s_mem_contents[14'h2bc8] = 8'h40;
s_mem_contents[14'h2bc9] = 8'h02;
s_mem_contents[14'h2bca] = 8'hd0;
s_mem_contents[14'h2bcb] = 8'hfe;
s_mem_contents[14'h2bcc] = 8'h68;
s_mem_contents[14'h2bcd] = 8'h49;
s_mem_contents[14'h2bce] = 8'h7d;
s_mem_contents[14'h2bcf] = 8'hdd;
s_mem_contents[14'h2bd0] = 8'h45;
s_mem_contents[14'h2bd1] = 8'h02;
s_mem_contents[14'h2bd2] = 8'hd0;
s_mem_contents[14'h2bd3] = 8'hfe;
s_mem_contents[14'h2bd4] = 8'hb5;
s_mem_contents[14'h2bd5] = 8'h02;
s_mem_contents[14'h2bd6] = 8'he8;
s_mem_contents[14'h2bd7] = 8'he0;
s_mem_contents[14'h2bd8] = 8'h02;
s_mem_contents[14'h2bd9] = 8'hd0;
s_mem_contents[14'h2bda] = 8'h02;
s_mem_contents[14'h2bdb] = 8'ha9;
s_mem_contents[14'h2bdc] = 8'hfe;
s_mem_contents[14'h2bdd] = 8'he0;
s_mem_contents[14'h2bde] = 8'h05;
s_mem_contents[14'h2bdf] = 8'hd0;
s_mem_contents[14'h2be0] = 8'hdb;
s_mem_contents[14'h2be1] = 8'hca;
s_mem_contents[14'h2be2] = 8'ha9;
s_mem_contents[14'h2be3] = 8'h02;
s_mem_contents[14'h2be4] = 8'h95;
s_mem_contents[14'h2be5] = 8'h02;
s_mem_contents[14'h2be6] = 8'ha9;
s_mem_contents[14'h2be7] = 8'hff;
s_mem_contents[14'h2be8] = 8'h48;
s_mem_contents[14'h2be9] = 8'h28;
s_mem_contents[14'h2bea] = 8'hd6;
s_mem_contents[14'h2beb] = 8'h02;
s_mem_contents[14'h2bec] = 8'h08;
s_mem_contents[14'h2bed] = 8'hb5;
s_mem_contents[14'h2bee] = 8'h02;
s_mem_contents[14'h2bef] = 8'hdd;
s_mem_contents[14'h2bf0] = 8'h40;
s_mem_contents[14'h2bf1] = 8'h02;
s_mem_contents[14'h2bf2] = 8'hd0;
s_mem_contents[14'h2bf3] = 8'hfe;
s_mem_contents[14'h2bf4] = 8'h68;
s_mem_contents[14'h2bf5] = 8'h49;
s_mem_contents[14'h2bf6] = 8'h7d;
s_mem_contents[14'h2bf7] = 8'hdd;
s_mem_contents[14'h2bf8] = 8'h45;
s_mem_contents[14'h2bf9] = 8'h02;
s_mem_contents[14'h2bfa] = 8'hd0;
s_mem_contents[14'h2bfb] = 8'hfe;
s_mem_contents[14'h2bfc] = 8'hb5;
s_mem_contents[14'h2bfd] = 8'h02;
s_mem_contents[14'h2bfe] = 8'hca;
s_mem_contents[14'h2bff] = 8'h30;
s_mem_contents[14'h2c00] = 8'h08;
s_mem_contents[14'h2c01] = 8'he0;
s_mem_contents[14'h2c02] = 8'h01;
s_mem_contents[14'h2c03] = 8'hd0;
s_mem_contents[14'h2c04] = 8'hdf;
s_mem_contents[14'h2c05] = 8'ha9;
s_mem_contents[14'h2c06] = 8'h81;
s_mem_contents[14'h2c07] = 8'hd0;
s_mem_contents[14'h2c08] = 8'hdb;
s_mem_contents[14'h2c09] = 8'had;
s_mem_contents[14'h2c0a] = 8'h00;
s_mem_contents[14'h2c0b] = 8'h02;
s_mem_contents[14'h2c0c] = 8'hc9;
s_mem_contents[14'h2c0d] = 8'h24;
s_mem_contents[14'h2c0e] = 8'hd0;
s_mem_contents[14'h2c0f] = 8'hfe;
s_mem_contents[14'h2c10] = 8'ha9;
s_mem_contents[14'h2c11] = 8'h25;
s_mem_contents[14'h2c12] = 8'h8d;
s_mem_contents[14'h2c13] = 8'h00;
s_mem_contents[14'h2c14] = 8'h02;
s_mem_contents[14'h2c15] = 8'ha2;
s_mem_contents[14'h2c16] = 8'h00;
s_mem_contents[14'h2c17] = 8'ha9;
s_mem_contents[14'h2c18] = 8'h7e;
s_mem_contents[14'h2c19] = 8'h9d;
s_mem_contents[14'h2c1a] = 8'h03;
s_mem_contents[14'h2c1b] = 8'h02;
s_mem_contents[14'h2c1c] = 8'ha9;
s_mem_contents[14'h2c1d] = 8'h00;
s_mem_contents[14'h2c1e] = 8'h48;
s_mem_contents[14'h2c1f] = 8'h28;
s_mem_contents[14'h2c20] = 8'hfe;
s_mem_contents[14'h2c21] = 8'h03;
s_mem_contents[14'h2c22] = 8'h02;
s_mem_contents[14'h2c23] = 8'h08;
s_mem_contents[14'h2c24] = 8'hbd;
s_mem_contents[14'h2c25] = 8'h03;
s_mem_contents[14'h2c26] = 8'h02;
s_mem_contents[14'h2c27] = 8'hdd;
s_mem_contents[14'h2c28] = 8'h40;
s_mem_contents[14'h2c29] = 8'h02;
s_mem_contents[14'h2c2a] = 8'hd0;
s_mem_contents[14'h2c2b] = 8'hfe;
s_mem_contents[14'h2c2c] = 8'h68;
s_mem_contents[14'h2c2d] = 8'h49;
s_mem_contents[14'h2c2e] = 8'h30;
s_mem_contents[14'h2c2f] = 8'hdd;
s_mem_contents[14'h2c30] = 8'h45;
s_mem_contents[14'h2c31] = 8'h02;
s_mem_contents[14'h2c32] = 8'hd0;
s_mem_contents[14'h2c33] = 8'hfe;
s_mem_contents[14'h2c34] = 8'hbd;
s_mem_contents[14'h2c35] = 8'h03;
s_mem_contents[14'h2c36] = 8'h02;
s_mem_contents[14'h2c37] = 8'he8;
s_mem_contents[14'h2c38] = 8'he0;
s_mem_contents[14'h2c39] = 8'h02;
s_mem_contents[14'h2c3a] = 8'hd0;
s_mem_contents[14'h2c3b] = 8'h02;
s_mem_contents[14'h2c3c] = 8'ha9;
s_mem_contents[14'h2c3d] = 8'hfe;
s_mem_contents[14'h2c3e] = 8'he0;
s_mem_contents[14'h2c3f] = 8'h05;
s_mem_contents[14'h2c40] = 8'hd0;
s_mem_contents[14'h2c41] = 8'hd7;
s_mem_contents[14'h2c42] = 8'hca;
s_mem_contents[14'h2c43] = 8'ha9;
s_mem_contents[14'h2c44] = 8'h02;
s_mem_contents[14'h2c45] = 8'h9d;
s_mem_contents[14'h2c46] = 8'h03;
s_mem_contents[14'h2c47] = 8'h02;
s_mem_contents[14'h2c48] = 8'ha9;
s_mem_contents[14'h2c49] = 8'h00;
s_mem_contents[14'h2c4a] = 8'h48;
s_mem_contents[14'h2c4b] = 8'h28;
s_mem_contents[14'h2c4c] = 8'hde;
s_mem_contents[14'h2c4d] = 8'h03;
s_mem_contents[14'h2c4e] = 8'h02;
s_mem_contents[14'h2c4f] = 8'h08;
s_mem_contents[14'h2c50] = 8'hbd;
s_mem_contents[14'h2c51] = 8'h03;
s_mem_contents[14'h2c52] = 8'h02;
s_mem_contents[14'h2c53] = 8'hdd;
s_mem_contents[14'h2c54] = 8'h40;
s_mem_contents[14'h2c55] = 8'h02;
s_mem_contents[14'h2c56] = 8'hd0;
s_mem_contents[14'h2c57] = 8'hfe;
s_mem_contents[14'h2c58] = 8'h68;
s_mem_contents[14'h2c59] = 8'h49;
s_mem_contents[14'h2c5a] = 8'h30;
s_mem_contents[14'h2c5b] = 8'hdd;
s_mem_contents[14'h2c5c] = 8'h45;
s_mem_contents[14'h2c5d] = 8'h02;
s_mem_contents[14'h2c5e] = 8'hd0;
s_mem_contents[14'h2c5f] = 8'hfe;
s_mem_contents[14'h2c60] = 8'hbd;
s_mem_contents[14'h2c61] = 8'h03;
s_mem_contents[14'h2c62] = 8'h02;
s_mem_contents[14'h2c63] = 8'hca;
s_mem_contents[14'h2c64] = 8'h30;
s_mem_contents[14'h2c65] = 8'h08;
s_mem_contents[14'h2c66] = 8'he0;
s_mem_contents[14'h2c67] = 8'h01;
s_mem_contents[14'h2c68] = 8'hd0;
s_mem_contents[14'h2c69] = 8'hdb;
s_mem_contents[14'h2c6a] = 8'ha9;
s_mem_contents[14'h2c6b] = 8'h81;
s_mem_contents[14'h2c6c] = 8'hd0;
s_mem_contents[14'h2c6d] = 8'hd7;
s_mem_contents[14'h2c6e] = 8'ha2;
s_mem_contents[14'h2c6f] = 8'h00;
s_mem_contents[14'h2c70] = 8'ha9;
s_mem_contents[14'h2c71] = 8'h7e;
s_mem_contents[14'h2c72] = 8'h9d;
s_mem_contents[14'h2c73] = 8'h03;
s_mem_contents[14'h2c74] = 8'h02;
s_mem_contents[14'h2c75] = 8'ha9;
s_mem_contents[14'h2c76] = 8'hff;
s_mem_contents[14'h2c77] = 8'h48;
s_mem_contents[14'h2c78] = 8'h28;
s_mem_contents[14'h2c79] = 8'hfe;
s_mem_contents[14'h2c7a] = 8'h03;
s_mem_contents[14'h2c7b] = 8'h02;
s_mem_contents[14'h2c7c] = 8'h08;
s_mem_contents[14'h2c7d] = 8'hbd;
s_mem_contents[14'h2c7e] = 8'h03;
s_mem_contents[14'h2c7f] = 8'h02;
s_mem_contents[14'h2c80] = 8'hdd;
s_mem_contents[14'h2c81] = 8'h40;
s_mem_contents[14'h2c82] = 8'h02;
s_mem_contents[14'h2c83] = 8'hd0;
s_mem_contents[14'h2c84] = 8'hfe;
s_mem_contents[14'h2c85] = 8'h68;
s_mem_contents[14'h2c86] = 8'h49;
s_mem_contents[14'h2c87] = 8'h7d;
s_mem_contents[14'h2c88] = 8'hdd;
s_mem_contents[14'h2c89] = 8'h45;
s_mem_contents[14'h2c8a] = 8'h02;
s_mem_contents[14'h2c8b] = 8'hd0;
s_mem_contents[14'h2c8c] = 8'hfe;
s_mem_contents[14'h2c8d] = 8'hbd;
s_mem_contents[14'h2c8e] = 8'h03;
s_mem_contents[14'h2c8f] = 8'h02;
s_mem_contents[14'h2c90] = 8'he8;
s_mem_contents[14'h2c91] = 8'he0;
s_mem_contents[14'h2c92] = 8'h02;
s_mem_contents[14'h2c93] = 8'hd0;
s_mem_contents[14'h2c94] = 8'h02;
s_mem_contents[14'h2c95] = 8'ha9;
s_mem_contents[14'h2c96] = 8'hfe;
s_mem_contents[14'h2c97] = 8'he0;
s_mem_contents[14'h2c98] = 8'h05;
s_mem_contents[14'h2c99] = 8'hd0;
s_mem_contents[14'h2c9a] = 8'hd7;
s_mem_contents[14'h2c9b] = 8'hca;
s_mem_contents[14'h2c9c] = 8'ha9;
s_mem_contents[14'h2c9d] = 8'h02;
s_mem_contents[14'h2c9e] = 8'h9d;
s_mem_contents[14'h2c9f] = 8'h03;
s_mem_contents[14'h2ca0] = 8'h02;
s_mem_contents[14'h2ca1] = 8'ha9;
s_mem_contents[14'h2ca2] = 8'hff;
s_mem_contents[14'h2ca3] = 8'h48;
s_mem_contents[14'h2ca4] = 8'h28;
s_mem_contents[14'h2ca5] = 8'hde;
s_mem_contents[14'h2ca6] = 8'h03;
s_mem_contents[14'h2ca7] = 8'h02;
s_mem_contents[14'h2ca8] = 8'h08;
s_mem_contents[14'h2ca9] = 8'hbd;
s_mem_contents[14'h2caa] = 8'h03;
s_mem_contents[14'h2cab] = 8'h02;
s_mem_contents[14'h2cac] = 8'hdd;
s_mem_contents[14'h2cad] = 8'h40;
s_mem_contents[14'h2cae] = 8'h02;
s_mem_contents[14'h2caf] = 8'hd0;
s_mem_contents[14'h2cb0] = 8'hfe;
s_mem_contents[14'h2cb1] = 8'h68;
s_mem_contents[14'h2cb2] = 8'h49;
s_mem_contents[14'h2cb3] = 8'h7d;
s_mem_contents[14'h2cb4] = 8'hdd;
s_mem_contents[14'h2cb5] = 8'h45;
s_mem_contents[14'h2cb6] = 8'h02;
s_mem_contents[14'h2cb7] = 8'hd0;
s_mem_contents[14'h2cb8] = 8'hfe;
s_mem_contents[14'h2cb9] = 8'hbd;
s_mem_contents[14'h2cba] = 8'h03;
s_mem_contents[14'h2cbb] = 8'h02;
s_mem_contents[14'h2cbc] = 8'hca;
s_mem_contents[14'h2cbd] = 8'h30;
s_mem_contents[14'h2cbe] = 8'h08;
s_mem_contents[14'h2cbf] = 8'he0;
s_mem_contents[14'h2cc0] = 8'h01;
s_mem_contents[14'h2cc1] = 8'hd0;
s_mem_contents[14'h2cc2] = 8'hdb;
s_mem_contents[14'h2cc3] = 8'ha9;
s_mem_contents[14'h2cc4] = 8'h81;
s_mem_contents[14'h2cc5] = 8'hd0;
s_mem_contents[14'h2cc6] = 8'hd7;
s_mem_contents[14'h2cc7] = 8'had;
s_mem_contents[14'h2cc8] = 8'h00;
s_mem_contents[14'h2cc9] = 8'h02;
s_mem_contents[14'h2cca] = 8'hc9;
s_mem_contents[14'h2ccb] = 8'h25;
s_mem_contents[14'h2ccc] = 8'hd0;
s_mem_contents[14'h2ccd] = 8'hfe;
s_mem_contents[14'h2cce] = 8'ha9;
s_mem_contents[14'h2ccf] = 8'h26;
s_mem_contents[14'h2cd0] = 8'h8d;
s_mem_contents[14'h2cd1] = 8'h00;
s_mem_contents[14'h2cd2] = 8'h02;
s_mem_contents[14'h2cd3] = 8'ha2;
s_mem_contents[14'h2cd4] = 8'h03;
s_mem_contents[14'h2cd5] = 8'hb5;
s_mem_contents[14'h2cd6] = 8'h12;
s_mem_contents[14'h2cd7] = 8'h8d;
s_mem_contents[14'h2cd8] = 8'h09;
s_mem_contents[14'h2cd9] = 8'h02;
s_mem_contents[14'h2cda] = 8'ha9;
s_mem_contents[14'h2cdb] = 8'h00;
s_mem_contents[14'h2cdc] = 8'h48;
s_mem_contents[14'h2cdd] = 8'hbd;
s_mem_contents[14'h2cde] = 8'h5a;
s_mem_contents[14'h2cdf] = 8'h02;
s_mem_contents[14'h2ce0] = 8'h28;
s_mem_contents[14'h2ce1] = 8'h20;
s_mem_contents[14'h2ce2] = 8'h08;
s_mem_contents[14'h2ce3] = 8'h02;
s_mem_contents[14'h2ce4] = 8'h08;
s_mem_contents[14'h2ce5] = 8'hdd;
s_mem_contents[14'h2ce6] = 8'h62;
s_mem_contents[14'h2ce7] = 8'h02;
s_mem_contents[14'h2ce8] = 8'hd0;
s_mem_contents[14'h2ce9] = 8'hfe;
s_mem_contents[14'h2cea] = 8'h68;
s_mem_contents[14'h2ceb] = 8'h49;
s_mem_contents[14'h2cec] = 8'h30;
s_mem_contents[14'h2ced] = 8'hdd;
s_mem_contents[14'h2cee] = 8'h66;
s_mem_contents[14'h2cef] = 8'h02;
s_mem_contents[14'h2cf0] = 8'hd0;
s_mem_contents[14'h2cf1] = 8'hfe;
s_mem_contents[14'h2cf2] = 8'hca;
s_mem_contents[14'h2cf3] = 8'h10;
s_mem_contents[14'h2cf4] = 8'he0;
s_mem_contents[14'h2cf5] = 8'ha2;
s_mem_contents[14'h2cf6] = 8'h03;
s_mem_contents[14'h2cf7] = 8'hb5;
s_mem_contents[14'h2cf8] = 8'h12;
s_mem_contents[14'h2cf9] = 8'h8d;
s_mem_contents[14'h2cfa] = 8'h09;
s_mem_contents[14'h2cfb] = 8'h02;
s_mem_contents[14'h2cfc] = 8'ha9;
s_mem_contents[14'h2cfd] = 8'hff;
s_mem_contents[14'h2cfe] = 8'h48;
s_mem_contents[14'h2cff] = 8'hbd;
s_mem_contents[14'h2d00] = 8'h5a;
s_mem_contents[14'h2d01] = 8'h02;
s_mem_contents[14'h2d02] = 8'h28;
s_mem_contents[14'h2d03] = 8'h20;
s_mem_contents[14'h2d04] = 8'h08;
s_mem_contents[14'h2d05] = 8'h02;
s_mem_contents[14'h2d06] = 8'h08;
s_mem_contents[14'h2d07] = 8'hdd;
s_mem_contents[14'h2d08] = 8'h62;
s_mem_contents[14'h2d09] = 8'h02;
s_mem_contents[14'h2d0a] = 8'hd0;
s_mem_contents[14'h2d0b] = 8'hfe;
s_mem_contents[14'h2d0c] = 8'h68;
s_mem_contents[14'h2d0d] = 8'h49;
s_mem_contents[14'h2d0e] = 8'h7d;
s_mem_contents[14'h2d0f] = 8'hdd;
s_mem_contents[14'h2d10] = 8'h66;
s_mem_contents[14'h2d11] = 8'h02;
s_mem_contents[14'h2d12] = 8'hd0;
s_mem_contents[14'h2d13] = 8'hfe;
s_mem_contents[14'h2d14] = 8'hca;
s_mem_contents[14'h2d15] = 8'h10;
s_mem_contents[14'h2d16] = 8'he0;
s_mem_contents[14'h2d17] = 8'ha2;
s_mem_contents[14'h2d18] = 8'h03;
s_mem_contents[14'h2d19] = 8'hb5;
s_mem_contents[14'h2d1a] = 8'h12;
s_mem_contents[14'h2d1b] = 8'h85;
s_mem_contents[14'h2d1c] = 8'h02;
s_mem_contents[14'h2d1d] = 8'ha9;
s_mem_contents[14'h2d1e] = 8'h00;
s_mem_contents[14'h2d1f] = 8'h48;
s_mem_contents[14'h2d20] = 8'hbd;
s_mem_contents[14'h2d21] = 8'h5a;
s_mem_contents[14'h2d22] = 8'h02;
s_mem_contents[14'h2d23] = 8'h28;
s_mem_contents[14'h2d24] = 8'h25;
s_mem_contents[14'h2d25] = 8'h02;
s_mem_contents[14'h2d26] = 8'h08;
s_mem_contents[14'h2d27] = 8'hdd;
s_mem_contents[14'h2d28] = 8'h62;
s_mem_contents[14'h2d29] = 8'h02;
s_mem_contents[14'h2d2a] = 8'hd0;
s_mem_contents[14'h2d2b] = 8'hfe;
s_mem_contents[14'h2d2c] = 8'h68;
s_mem_contents[14'h2d2d] = 8'h49;
s_mem_contents[14'h2d2e] = 8'h30;
s_mem_contents[14'h2d2f] = 8'hdd;
s_mem_contents[14'h2d30] = 8'h66;
s_mem_contents[14'h2d31] = 8'h02;
s_mem_contents[14'h2d32] = 8'hd0;
s_mem_contents[14'h2d33] = 8'hfe;
s_mem_contents[14'h2d34] = 8'hca;
s_mem_contents[14'h2d35] = 8'h10;
s_mem_contents[14'h2d36] = 8'he2;
s_mem_contents[14'h2d37] = 8'ha2;
s_mem_contents[14'h2d38] = 8'h03;
s_mem_contents[14'h2d39] = 8'hb5;
s_mem_contents[14'h2d3a] = 8'h12;
s_mem_contents[14'h2d3b] = 8'h85;
s_mem_contents[14'h2d3c] = 8'h02;
s_mem_contents[14'h2d3d] = 8'ha9;
s_mem_contents[14'h2d3e] = 8'hff;
s_mem_contents[14'h2d3f] = 8'h48;
s_mem_contents[14'h2d40] = 8'hbd;
s_mem_contents[14'h2d41] = 8'h5a;
s_mem_contents[14'h2d42] = 8'h02;
s_mem_contents[14'h2d43] = 8'h28;
s_mem_contents[14'h2d44] = 8'h25;
s_mem_contents[14'h2d45] = 8'h02;
s_mem_contents[14'h2d46] = 8'h08;
s_mem_contents[14'h2d47] = 8'hdd;
s_mem_contents[14'h2d48] = 8'h62;
s_mem_contents[14'h2d49] = 8'h02;
s_mem_contents[14'h2d4a] = 8'hd0;
s_mem_contents[14'h2d4b] = 8'hfe;
s_mem_contents[14'h2d4c] = 8'h68;
s_mem_contents[14'h2d4d] = 8'h49;
s_mem_contents[14'h2d4e] = 8'h7d;
s_mem_contents[14'h2d4f] = 8'hdd;
s_mem_contents[14'h2d50] = 8'h66;
s_mem_contents[14'h2d51] = 8'h02;
s_mem_contents[14'h2d52] = 8'hd0;
s_mem_contents[14'h2d53] = 8'hfe;
s_mem_contents[14'h2d54] = 8'hca;
s_mem_contents[14'h2d55] = 8'h10;
s_mem_contents[14'h2d56] = 8'he2;
s_mem_contents[14'h2d57] = 8'ha2;
s_mem_contents[14'h2d58] = 8'h03;
s_mem_contents[14'h2d59] = 8'hb5;
s_mem_contents[14'h2d5a] = 8'h12;
s_mem_contents[14'h2d5b] = 8'h8d;
s_mem_contents[14'h2d5c] = 8'h03;
s_mem_contents[14'h2d5d] = 8'h02;
s_mem_contents[14'h2d5e] = 8'ha9;
s_mem_contents[14'h2d5f] = 8'h00;
s_mem_contents[14'h2d60] = 8'h48;
s_mem_contents[14'h2d61] = 8'hbd;
s_mem_contents[14'h2d62] = 8'h5a;
s_mem_contents[14'h2d63] = 8'h02;
s_mem_contents[14'h2d64] = 8'h28;
s_mem_contents[14'h2d65] = 8'h2d;
s_mem_contents[14'h2d66] = 8'h03;
s_mem_contents[14'h2d67] = 8'h02;
s_mem_contents[14'h2d68] = 8'h08;
s_mem_contents[14'h2d69] = 8'hdd;
s_mem_contents[14'h2d6a] = 8'h62;
s_mem_contents[14'h2d6b] = 8'h02;
s_mem_contents[14'h2d6c] = 8'hd0;
s_mem_contents[14'h2d6d] = 8'hfe;
s_mem_contents[14'h2d6e] = 8'h68;
s_mem_contents[14'h2d6f] = 8'h49;
s_mem_contents[14'h2d70] = 8'h30;
s_mem_contents[14'h2d71] = 8'hdd;
s_mem_contents[14'h2d72] = 8'h66;
s_mem_contents[14'h2d73] = 8'h02;
s_mem_contents[14'h2d74] = 8'hd0;
s_mem_contents[14'h2d75] = 8'hfe;
s_mem_contents[14'h2d76] = 8'hca;
s_mem_contents[14'h2d77] = 8'h10;
s_mem_contents[14'h2d78] = 8'he0;
s_mem_contents[14'h2d79] = 8'ha2;
s_mem_contents[14'h2d7a] = 8'h03;
s_mem_contents[14'h2d7b] = 8'hb5;
s_mem_contents[14'h2d7c] = 8'h12;
s_mem_contents[14'h2d7d] = 8'h8d;
s_mem_contents[14'h2d7e] = 8'h03;
s_mem_contents[14'h2d7f] = 8'h02;
s_mem_contents[14'h2d80] = 8'ha9;
s_mem_contents[14'h2d81] = 8'hff;
s_mem_contents[14'h2d82] = 8'h48;
s_mem_contents[14'h2d83] = 8'hbd;
s_mem_contents[14'h2d84] = 8'h5a;
s_mem_contents[14'h2d85] = 8'h02;
s_mem_contents[14'h2d86] = 8'h28;
s_mem_contents[14'h2d87] = 8'h2d;
s_mem_contents[14'h2d88] = 8'h03;
s_mem_contents[14'h2d89] = 8'h02;
s_mem_contents[14'h2d8a] = 8'h08;
s_mem_contents[14'h2d8b] = 8'hdd;
s_mem_contents[14'h2d8c] = 8'h62;
s_mem_contents[14'h2d8d] = 8'h02;
s_mem_contents[14'h2d8e] = 8'hd0;
s_mem_contents[14'h2d8f] = 8'hfe;
s_mem_contents[14'h2d90] = 8'h68;
s_mem_contents[14'h2d91] = 8'h49;
s_mem_contents[14'h2d92] = 8'h7d;
s_mem_contents[14'h2d93] = 8'hdd;
s_mem_contents[14'h2d94] = 8'h66;
s_mem_contents[14'h2d95] = 8'h02;
s_mem_contents[14'h2d96] = 8'hd0;
s_mem_contents[14'h2d97] = 8'hfe;
s_mem_contents[14'h2d98] = 8'hca;
s_mem_contents[14'h2d99] = 8'h10;
s_mem_contents[14'h2d9a] = 8'h02;
s_mem_contents[14'h2d9b] = 8'ha2;
s_mem_contents[14'h2d9c] = 8'h03;
s_mem_contents[14'h2d9d] = 8'ha9;
s_mem_contents[14'h2d9e] = 8'h00;
s_mem_contents[14'h2d9f] = 8'h48;
s_mem_contents[14'h2da0] = 8'hbd;
s_mem_contents[14'h2da1] = 8'h5a;
s_mem_contents[14'h2da2] = 8'h02;
s_mem_contents[14'h2da3] = 8'h28;
s_mem_contents[14'h2da4] = 8'h35;
s_mem_contents[14'h2da5] = 8'h12;
s_mem_contents[14'h2da6] = 8'h08;
s_mem_contents[14'h2da7] = 8'hdd;
s_mem_contents[14'h2da8] = 8'h62;
s_mem_contents[14'h2da9] = 8'h02;
s_mem_contents[14'h2daa] = 8'hd0;
s_mem_contents[14'h2dab] = 8'hfe;
s_mem_contents[14'h2dac] = 8'h68;
s_mem_contents[14'h2dad] = 8'h49;
s_mem_contents[14'h2dae] = 8'h30;
s_mem_contents[14'h2daf] = 8'hdd;
s_mem_contents[14'h2db0] = 8'h66;
s_mem_contents[14'h2db1] = 8'h02;
s_mem_contents[14'h2db2] = 8'hd0;
s_mem_contents[14'h2db3] = 8'hfe;
s_mem_contents[14'h2db4] = 8'hca;
s_mem_contents[14'h2db5] = 8'h10;
s_mem_contents[14'h2db6] = 8'he6;
s_mem_contents[14'h2db7] = 8'ha2;
s_mem_contents[14'h2db8] = 8'h03;
s_mem_contents[14'h2db9] = 8'ha9;
s_mem_contents[14'h2dba] = 8'hff;
s_mem_contents[14'h2dbb] = 8'h48;
s_mem_contents[14'h2dbc] = 8'hbd;
s_mem_contents[14'h2dbd] = 8'h5a;
s_mem_contents[14'h2dbe] = 8'h02;
s_mem_contents[14'h2dbf] = 8'h28;
s_mem_contents[14'h2dc0] = 8'h35;
s_mem_contents[14'h2dc1] = 8'h12;
s_mem_contents[14'h2dc2] = 8'h08;
s_mem_contents[14'h2dc3] = 8'hdd;
s_mem_contents[14'h2dc4] = 8'h62;
s_mem_contents[14'h2dc5] = 8'h02;
s_mem_contents[14'h2dc6] = 8'hd0;
s_mem_contents[14'h2dc7] = 8'hfe;
s_mem_contents[14'h2dc8] = 8'h68;
s_mem_contents[14'h2dc9] = 8'h49;
s_mem_contents[14'h2dca] = 8'h7d;
s_mem_contents[14'h2dcb] = 8'hdd;
s_mem_contents[14'h2dcc] = 8'h66;
s_mem_contents[14'h2dcd] = 8'h02;
s_mem_contents[14'h2dce] = 8'hd0;
s_mem_contents[14'h2dcf] = 8'hfe;
s_mem_contents[14'h2dd0] = 8'hca;
s_mem_contents[14'h2dd1] = 8'h10;
s_mem_contents[14'h2dd2] = 8'he6;
s_mem_contents[14'h2dd3] = 8'ha2;
s_mem_contents[14'h2dd4] = 8'h03;
s_mem_contents[14'h2dd5] = 8'ha9;
s_mem_contents[14'h2dd6] = 8'h00;
s_mem_contents[14'h2dd7] = 8'h48;
s_mem_contents[14'h2dd8] = 8'hbd;
s_mem_contents[14'h2dd9] = 8'h5a;
s_mem_contents[14'h2dda] = 8'h02;
s_mem_contents[14'h2ddb] = 8'h28;
s_mem_contents[14'h2ddc] = 8'h3d;
s_mem_contents[14'h2ddd] = 8'h4e;
s_mem_contents[14'h2dde] = 8'h02;
s_mem_contents[14'h2ddf] = 8'h08;
s_mem_contents[14'h2de0] = 8'hdd;
s_mem_contents[14'h2de1] = 8'h62;
s_mem_contents[14'h2de2] = 8'h02;
s_mem_contents[14'h2de3] = 8'hd0;
s_mem_contents[14'h2de4] = 8'hfe;
s_mem_contents[14'h2de5] = 8'h68;
s_mem_contents[14'h2de6] = 8'h49;
s_mem_contents[14'h2de7] = 8'h30;
s_mem_contents[14'h2de8] = 8'hdd;
s_mem_contents[14'h2de9] = 8'h66;
s_mem_contents[14'h2dea] = 8'h02;
s_mem_contents[14'h2deb] = 8'hd0;
s_mem_contents[14'h2dec] = 8'hfe;
s_mem_contents[14'h2ded] = 8'hca;
s_mem_contents[14'h2dee] = 8'h10;
s_mem_contents[14'h2def] = 8'he5;
s_mem_contents[14'h2df0] = 8'ha2;
s_mem_contents[14'h2df1] = 8'h03;
s_mem_contents[14'h2df2] = 8'ha9;
s_mem_contents[14'h2df3] = 8'hff;
s_mem_contents[14'h2df4] = 8'h48;
s_mem_contents[14'h2df5] = 8'hbd;
s_mem_contents[14'h2df6] = 8'h5a;
s_mem_contents[14'h2df7] = 8'h02;
s_mem_contents[14'h2df8] = 8'h28;
s_mem_contents[14'h2df9] = 8'h3d;
s_mem_contents[14'h2dfa] = 8'h4e;
s_mem_contents[14'h2dfb] = 8'h02;
s_mem_contents[14'h2dfc] = 8'h08;
s_mem_contents[14'h2dfd] = 8'hdd;
s_mem_contents[14'h2dfe] = 8'h62;
s_mem_contents[14'h2dff] = 8'h02;
s_mem_contents[14'h2e00] = 8'hd0;
s_mem_contents[14'h2e01] = 8'hfe;
s_mem_contents[14'h2e02] = 8'h68;
s_mem_contents[14'h2e03] = 8'h49;
s_mem_contents[14'h2e04] = 8'h7d;
s_mem_contents[14'h2e05] = 8'hdd;
s_mem_contents[14'h2e06] = 8'h66;
s_mem_contents[14'h2e07] = 8'h02;
s_mem_contents[14'h2e08] = 8'hd0;
s_mem_contents[14'h2e09] = 8'hfe;
s_mem_contents[14'h2e0a] = 8'hca;
s_mem_contents[14'h2e0b] = 8'h10;
s_mem_contents[14'h2e0c] = 8'he5;
s_mem_contents[14'h2e0d] = 8'ha0;
s_mem_contents[14'h2e0e] = 8'h03;
s_mem_contents[14'h2e0f] = 8'ha9;
s_mem_contents[14'h2e10] = 8'h00;
s_mem_contents[14'h2e11] = 8'h48;
s_mem_contents[14'h2e12] = 8'hb9;
s_mem_contents[14'h2e13] = 8'h5a;
s_mem_contents[14'h2e14] = 8'h02;
s_mem_contents[14'h2e15] = 8'h28;
s_mem_contents[14'h2e16] = 8'h39;
s_mem_contents[14'h2e17] = 8'h4e;
s_mem_contents[14'h2e18] = 8'h02;
s_mem_contents[14'h2e19] = 8'h08;
s_mem_contents[14'h2e1a] = 8'hd9;
s_mem_contents[14'h2e1b] = 8'h62;
s_mem_contents[14'h2e1c] = 8'h02;
s_mem_contents[14'h2e1d] = 8'hd0;
s_mem_contents[14'h2e1e] = 8'hfe;
s_mem_contents[14'h2e1f] = 8'h68;
s_mem_contents[14'h2e20] = 8'h49;
s_mem_contents[14'h2e21] = 8'h30;
s_mem_contents[14'h2e22] = 8'hd9;
s_mem_contents[14'h2e23] = 8'h66;
s_mem_contents[14'h2e24] = 8'h02;
s_mem_contents[14'h2e25] = 8'hd0;
s_mem_contents[14'h2e26] = 8'hfe;
s_mem_contents[14'h2e27] = 8'h88;
s_mem_contents[14'h2e28] = 8'h10;
s_mem_contents[14'h2e29] = 8'he5;
s_mem_contents[14'h2e2a] = 8'ha0;
s_mem_contents[14'h2e2b] = 8'h03;
s_mem_contents[14'h2e2c] = 8'ha9;
s_mem_contents[14'h2e2d] = 8'hff;
s_mem_contents[14'h2e2e] = 8'h48;
s_mem_contents[14'h2e2f] = 8'hb9;
s_mem_contents[14'h2e30] = 8'h5a;
s_mem_contents[14'h2e31] = 8'h02;
s_mem_contents[14'h2e32] = 8'h28;
s_mem_contents[14'h2e33] = 8'h39;
s_mem_contents[14'h2e34] = 8'h4e;
s_mem_contents[14'h2e35] = 8'h02;
s_mem_contents[14'h2e36] = 8'h08;
s_mem_contents[14'h2e37] = 8'hd9;
s_mem_contents[14'h2e38] = 8'h62;
s_mem_contents[14'h2e39] = 8'h02;
s_mem_contents[14'h2e3a] = 8'hd0;
s_mem_contents[14'h2e3b] = 8'hfe;
s_mem_contents[14'h2e3c] = 8'h68;
s_mem_contents[14'h2e3d] = 8'h49;
s_mem_contents[14'h2e3e] = 8'h7d;
s_mem_contents[14'h2e3f] = 8'hd9;
s_mem_contents[14'h2e40] = 8'h66;
s_mem_contents[14'h2e41] = 8'h02;
s_mem_contents[14'h2e42] = 8'hd0;
s_mem_contents[14'h2e43] = 8'hfe;
s_mem_contents[14'h2e44] = 8'h88;
s_mem_contents[14'h2e45] = 8'h10;
s_mem_contents[14'h2e46] = 8'he5;
s_mem_contents[14'h2e47] = 8'ha2;
s_mem_contents[14'h2e48] = 8'h06;
s_mem_contents[14'h2e49] = 8'ha0;
s_mem_contents[14'h2e4a] = 8'h03;
s_mem_contents[14'h2e4b] = 8'ha9;
s_mem_contents[14'h2e4c] = 8'h00;
s_mem_contents[14'h2e4d] = 8'h48;
s_mem_contents[14'h2e4e] = 8'hb9;
s_mem_contents[14'h2e4f] = 8'h5a;
s_mem_contents[14'h2e50] = 8'h02;
s_mem_contents[14'h2e51] = 8'h28;
s_mem_contents[14'h2e52] = 8'h21;
s_mem_contents[14'h2e53] = 8'h30;
s_mem_contents[14'h2e54] = 8'h08;
s_mem_contents[14'h2e55] = 8'hd9;
s_mem_contents[14'h2e56] = 8'h62;
s_mem_contents[14'h2e57] = 8'h02;
s_mem_contents[14'h2e58] = 8'hd0;
s_mem_contents[14'h2e59] = 8'hfe;
s_mem_contents[14'h2e5a] = 8'h68;
s_mem_contents[14'h2e5b] = 8'h49;
s_mem_contents[14'h2e5c] = 8'h30;
s_mem_contents[14'h2e5d] = 8'hd9;
s_mem_contents[14'h2e5e] = 8'h66;
s_mem_contents[14'h2e5f] = 8'h02;
s_mem_contents[14'h2e60] = 8'hd0;
s_mem_contents[14'h2e61] = 8'hfe;
s_mem_contents[14'h2e62] = 8'hca;
s_mem_contents[14'h2e63] = 8'hca;
s_mem_contents[14'h2e64] = 8'h88;
s_mem_contents[14'h2e65] = 8'h10;
s_mem_contents[14'h2e66] = 8'he4;
s_mem_contents[14'h2e67] = 8'ha2;
s_mem_contents[14'h2e68] = 8'h06;
s_mem_contents[14'h2e69] = 8'ha0;
s_mem_contents[14'h2e6a] = 8'h03;
s_mem_contents[14'h2e6b] = 8'ha9;
s_mem_contents[14'h2e6c] = 8'hff;
s_mem_contents[14'h2e6d] = 8'h48;
s_mem_contents[14'h2e6e] = 8'hb9;
s_mem_contents[14'h2e6f] = 8'h5a;
s_mem_contents[14'h2e70] = 8'h02;
s_mem_contents[14'h2e71] = 8'h28;
s_mem_contents[14'h2e72] = 8'h21;
s_mem_contents[14'h2e73] = 8'h30;
s_mem_contents[14'h2e74] = 8'h08;
s_mem_contents[14'h2e75] = 8'hd9;
s_mem_contents[14'h2e76] = 8'h62;
s_mem_contents[14'h2e77] = 8'h02;
s_mem_contents[14'h2e78] = 8'hd0;
s_mem_contents[14'h2e79] = 8'hfe;
s_mem_contents[14'h2e7a] = 8'h68;
s_mem_contents[14'h2e7b] = 8'h49;
s_mem_contents[14'h2e7c] = 8'h7d;
s_mem_contents[14'h2e7d] = 8'hd9;
s_mem_contents[14'h2e7e] = 8'h66;
s_mem_contents[14'h2e7f] = 8'h02;
s_mem_contents[14'h2e80] = 8'hd0;
s_mem_contents[14'h2e81] = 8'hfe;
s_mem_contents[14'h2e82] = 8'hca;
s_mem_contents[14'h2e83] = 8'hca;
s_mem_contents[14'h2e84] = 8'h88;
s_mem_contents[14'h2e85] = 8'h10;
s_mem_contents[14'h2e86] = 8'he4;
s_mem_contents[14'h2e87] = 8'ha0;
s_mem_contents[14'h2e88] = 8'h03;
s_mem_contents[14'h2e89] = 8'ha9;
s_mem_contents[14'h2e8a] = 8'h00;
s_mem_contents[14'h2e8b] = 8'h48;
s_mem_contents[14'h2e8c] = 8'hb9;
s_mem_contents[14'h2e8d] = 8'h5a;
s_mem_contents[14'h2e8e] = 8'h02;
s_mem_contents[14'h2e8f] = 8'h28;
s_mem_contents[14'h2e90] = 8'h31;
s_mem_contents[14'h2e91] = 8'h30;
s_mem_contents[14'h2e92] = 8'h08;
s_mem_contents[14'h2e93] = 8'hd9;
s_mem_contents[14'h2e94] = 8'h62;
s_mem_contents[14'h2e95] = 8'h02;
s_mem_contents[14'h2e96] = 8'hd0;
s_mem_contents[14'h2e97] = 8'hfe;
s_mem_contents[14'h2e98] = 8'h68;
s_mem_contents[14'h2e99] = 8'h49;
s_mem_contents[14'h2e9a] = 8'h30;
s_mem_contents[14'h2e9b] = 8'hd9;
s_mem_contents[14'h2e9c] = 8'h66;
s_mem_contents[14'h2e9d] = 8'h02;
s_mem_contents[14'h2e9e] = 8'hd0;
s_mem_contents[14'h2e9f] = 8'hfe;
s_mem_contents[14'h2ea0] = 8'h88;
s_mem_contents[14'h2ea1] = 8'h10;
s_mem_contents[14'h2ea2] = 8'he6;
s_mem_contents[14'h2ea3] = 8'ha0;
s_mem_contents[14'h2ea4] = 8'h03;
s_mem_contents[14'h2ea5] = 8'ha9;
s_mem_contents[14'h2ea6] = 8'hff;
s_mem_contents[14'h2ea7] = 8'h48;
s_mem_contents[14'h2ea8] = 8'hb9;
s_mem_contents[14'h2ea9] = 8'h5a;
s_mem_contents[14'h2eaa] = 8'h02;
s_mem_contents[14'h2eab] = 8'h28;
s_mem_contents[14'h2eac] = 8'h31;
s_mem_contents[14'h2ead] = 8'h30;
s_mem_contents[14'h2eae] = 8'h08;
s_mem_contents[14'h2eaf] = 8'hd9;
s_mem_contents[14'h2eb0] = 8'h62;
s_mem_contents[14'h2eb1] = 8'h02;
s_mem_contents[14'h2eb2] = 8'hd0;
s_mem_contents[14'h2eb3] = 8'hfe;
s_mem_contents[14'h2eb4] = 8'h68;
s_mem_contents[14'h2eb5] = 8'h49;
s_mem_contents[14'h2eb6] = 8'h7d;
s_mem_contents[14'h2eb7] = 8'hd9;
s_mem_contents[14'h2eb8] = 8'h66;
s_mem_contents[14'h2eb9] = 8'h02;
s_mem_contents[14'h2eba] = 8'hd0;
s_mem_contents[14'h2ebb] = 8'hfe;
s_mem_contents[14'h2ebc] = 8'h88;
s_mem_contents[14'h2ebd] = 8'h10;
s_mem_contents[14'h2ebe] = 8'he6;
s_mem_contents[14'h2ebf] = 8'had;
s_mem_contents[14'h2ec0] = 8'h00;
s_mem_contents[14'h2ec1] = 8'h02;
s_mem_contents[14'h2ec2] = 8'hc9;
s_mem_contents[14'h2ec3] = 8'h26;
s_mem_contents[14'h2ec4] = 8'hd0;
s_mem_contents[14'h2ec5] = 8'hfe;
s_mem_contents[14'h2ec6] = 8'ha9;
s_mem_contents[14'h2ec7] = 8'h27;
s_mem_contents[14'h2ec8] = 8'h8d;
s_mem_contents[14'h2ec9] = 8'h00;
s_mem_contents[14'h2eca] = 8'h02;
s_mem_contents[14'h2ecb] = 8'ha2;
s_mem_contents[14'h2ecc] = 8'h03;
s_mem_contents[14'h2ecd] = 8'hb5;
s_mem_contents[14'h2ece] = 8'h16;
s_mem_contents[14'h2ecf] = 8'h8d;
s_mem_contents[14'h2ed0] = 8'h0c;
s_mem_contents[14'h2ed1] = 8'h02;
s_mem_contents[14'h2ed2] = 8'ha9;
s_mem_contents[14'h2ed3] = 8'h00;
s_mem_contents[14'h2ed4] = 8'h48;
s_mem_contents[14'h2ed5] = 8'hbd;
s_mem_contents[14'h2ed6] = 8'h5e;
s_mem_contents[14'h2ed7] = 8'h02;
s_mem_contents[14'h2ed8] = 8'h28;
s_mem_contents[14'h2ed9] = 8'h20;
s_mem_contents[14'h2eda] = 8'h0b;
s_mem_contents[14'h2edb] = 8'h02;
s_mem_contents[14'h2edc] = 8'h08;
s_mem_contents[14'h2edd] = 8'hdd;
s_mem_contents[14'h2ede] = 8'h62;
s_mem_contents[14'h2edf] = 8'h02;
s_mem_contents[14'h2ee0] = 8'hd0;
s_mem_contents[14'h2ee1] = 8'hfe;
s_mem_contents[14'h2ee2] = 8'h68;
s_mem_contents[14'h2ee3] = 8'h49;
s_mem_contents[14'h2ee4] = 8'h30;
s_mem_contents[14'h2ee5] = 8'hdd;
s_mem_contents[14'h2ee6] = 8'h66;
s_mem_contents[14'h2ee7] = 8'h02;
s_mem_contents[14'h2ee8] = 8'hd0;
s_mem_contents[14'h2ee9] = 8'hfe;
s_mem_contents[14'h2eea] = 8'hca;
s_mem_contents[14'h2eeb] = 8'h10;
s_mem_contents[14'h2eec] = 8'he0;
s_mem_contents[14'h2eed] = 8'ha2;
s_mem_contents[14'h2eee] = 8'h03;
s_mem_contents[14'h2eef] = 8'hb5;
s_mem_contents[14'h2ef0] = 8'h16;
s_mem_contents[14'h2ef1] = 8'h8d;
s_mem_contents[14'h2ef2] = 8'h0c;
s_mem_contents[14'h2ef3] = 8'h02;
s_mem_contents[14'h2ef4] = 8'ha9;
s_mem_contents[14'h2ef5] = 8'hff;
s_mem_contents[14'h2ef6] = 8'h48;
s_mem_contents[14'h2ef7] = 8'hbd;
s_mem_contents[14'h2ef8] = 8'h5e;
s_mem_contents[14'h2ef9] = 8'h02;
s_mem_contents[14'h2efa] = 8'h28;
s_mem_contents[14'h2efb] = 8'h20;
s_mem_contents[14'h2efc] = 8'h0b;
s_mem_contents[14'h2efd] = 8'h02;
s_mem_contents[14'h2efe] = 8'h08;
s_mem_contents[14'h2eff] = 8'hdd;
s_mem_contents[14'h2f00] = 8'h62;
s_mem_contents[14'h2f01] = 8'h02;
s_mem_contents[14'h2f02] = 8'hd0;
s_mem_contents[14'h2f03] = 8'hfe;
s_mem_contents[14'h2f04] = 8'h68;
s_mem_contents[14'h2f05] = 8'h49;
s_mem_contents[14'h2f06] = 8'h7d;
s_mem_contents[14'h2f07] = 8'hdd;
s_mem_contents[14'h2f08] = 8'h66;
s_mem_contents[14'h2f09] = 8'h02;
s_mem_contents[14'h2f0a] = 8'hd0;
s_mem_contents[14'h2f0b] = 8'hfe;
s_mem_contents[14'h2f0c] = 8'hca;
s_mem_contents[14'h2f0d] = 8'h10;
s_mem_contents[14'h2f0e] = 8'he0;
s_mem_contents[14'h2f0f] = 8'ha2;
s_mem_contents[14'h2f10] = 8'h03;
s_mem_contents[14'h2f11] = 8'hb5;
s_mem_contents[14'h2f12] = 8'h16;
s_mem_contents[14'h2f13] = 8'h85;
s_mem_contents[14'h2f14] = 8'h02;
s_mem_contents[14'h2f15] = 8'ha9;
s_mem_contents[14'h2f16] = 8'h00;
s_mem_contents[14'h2f17] = 8'h48;
s_mem_contents[14'h2f18] = 8'hbd;
s_mem_contents[14'h2f19] = 8'h5e;
s_mem_contents[14'h2f1a] = 8'h02;
s_mem_contents[14'h2f1b] = 8'h28;
s_mem_contents[14'h2f1c] = 8'h45;
s_mem_contents[14'h2f1d] = 8'h02;
s_mem_contents[14'h2f1e] = 8'h08;
s_mem_contents[14'h2f1f] = 8'hdd;
s_mem_contents[14'h2f20] = 8'h62;
s_mem_contents[14'h2f21] = 8'h02;
s_mem_contents[14'h2f22] = 8'hd0;
s_mem_contents[14'h2f23] = 8'hfe;
s_mem_contents[14'h2f24] = 8'h68;
s_mem_contents[14'h2f25] = 8'h49;
s_mem_contents[14'h2f26] = 8'h30;
s_mem_contents[14'h2f27] = 8'hdd;
s_mem_contents[14'h2f28] = 8'h66;
s_mem_contents[14'h2f29] = 8'h02;
s_mem_contents[14'h2f2a] = 8'hd0;
s_mem_contents[14'h2f2b] = 8'hfe;
s_mem_contents[14'h2f2c] = 8'hca;
s_mem_contents[14'h2f2d] = 8'h10;
s_mem_contents[14'h2f2e] = 8'he2;
s_mem_contents[14'h2f2f] = 8'ha2;
s_mem_contents[14'h2f30] = 8'h03;
s_mem_contents[14'h2f31] = 8'hb5;
s_mem_contents[14'h2f32] = 8'h16;
s_mem_contents[14'h2f33] = 8'h85;
s_mem_contents[14'h2f34] = 8'h02;
s_mem_contents[14'h2f35] = 8'ha9;
s_mem_contents[14'h2f36] = 8'hff;
s_mem_contents[14'h2f37] = 8'h48;
s_mem_contents[14'h2f38] = 8'hbd;
s_mem_contents[14'h2f39] = 8'h5e;
s_mem_contents[14'h2f3a] = 8'h02;
s_mem_contents[14'h2f3b] = 8'h28;
s_mem_contents[14'h2f3c] = 8'h45;
s_mem_contents[14'h2f3d] = 8'h02;
s_mem_contents[14'h2f3e] = 8'h08;
s_mem_contents[14'h2f3f] = 8'hdd;
s_mem_contents[14'h2f40] = 8'h62;
s_mem_contents[14'h2f41] = 8'h02;
s_mem_contents[14'h2f42] = 8'hd0;
s_mem_contents[14'h2f43] = 8'hfe;
s_mem_contents[14'h2f44] = 8'h68;
s_mem_contents[14'h2f45] = 8'h49;
s_mem_contents[14'h2f46] = 8'h7d;
s_mem_contents[14'h2f47] = 8'hdd;
s_mem_contents[14'h2f48] = 8'h66;
s_mem_contents[14'h2f49] = 8'h02;
s_mem_contents[14'h2f4a] = 8'hd0;
s_mem_contents[14'h2f4b] = 8'hfe;
s_mem_contents[14'h2f4c] = 8'hca;
s_mem_contents[14'h2f4d] = 8'h10;
s_mem_contents[14'h2f4e] = 8'he2;
s_mem_contents[14'h2f4f] = 8'ha2;
s_mem_contents[14'h2f50] = 8'h03;
s_mem_contents[14'h2f51] = 8'hb5;
s_mem_contents[14'h2f52] = 8'h16;
s_mem_contents[14'h2f53] = 8'h8d;
s_mem_contents[14'h2f54] = 8'h03;
s_mem_contents[14'h2f55] = 8'h02;
s_mem_contents[14'h2f56] = 8'ha9;
s_mem_contents[14'h2f57] = 8'h00;
s_mem_contents[14'h2f58] = 8'h48;
s_mem_contents[14'h2f59] = 8'hbd;
s_mem_contents[14'h2f5a] = 8'h5e;
s_mem_contents[14'h2f5b] = 8'h02;
s_mem_contents[14'h2f5c] = 8'h28;
s_mem_contents[14'h2f5d] = 8'h4d;
s_mem_contents[14'h2f5e] = 8'h03;
s_mem_contents[14'h2f5f] = 8'h02;
s_mem_contents[14'h2f60] = 8'h08;
s_mem_contents[14'h2f61] = 8'hdd;
s_mem_contents[14'h2f62] = 8'h62;
s_mem_contents[14'h2f63] = 8'h02;
s_mem_contents[14'h2f64] = 8'hd0;
s_mem_contents[14'h2f65] = 8'hfe;
s_mem_contents[14'h2f66] = 8'h68;
s_mem_contents[14'h2f67] = 8'h49;
s_mem_contents[14'h2f68] = 8'h30;
s_mem_contents[14'h2f69] = 8'hdd;
s_mem_contents[14'h2f6a] = 8'h66;
s_mem_contents[14'h2f6b] = 8'h02;
s_mem_contents[14'h2f6c] = 8'hd0;
s_mem_contents[14'h2f6d] = 8'hfe;
s_mem_contents[14'h2f6e] = 8'hca;
s_mem_contents[14'h2f6f] = 8'h10;
s_mem_contents[14'h2f70] = 8'he0;
s_mem_contents[14'h2f71] = 8'ha2;
s_mem_contents[14'h2f72] = 8'h03;
s_mem_contents[14'h2f73] = 8'hb5;
s_mem_contents[14'h2f74] = 8'h16;
s_mem_contents[14'h2f75] = 8'h8d;
s_mem_contents[14'h2f76] = 8'h03;
s_mem_contents[14'h2f77] = 8'h02;
s_mem_contents[14'h2f78] = 8'ha9;
s_mem_contents[14'h2f79] = 8'hff;
s_mem_contents[14'h2f7a] = 8'h48;
s_mem_contents[14'h2f7b] = 8'hbd;
s_mem_contents[14'h2f7c] = 8'h5e;
s_mem_contents[14'h2f7d] = 8'h02;
s_mem_contents[14'h2f7e] = 8'h28;
s_mem_contents[14'h2f7f] = 8'h4d;
s_mem_contents[14'h2f80] = 8'h03;
s_mem_contents[14'h2f81] = 8'h02;
s_mem_contents[14'h2f82] = 8'h08;
s_mem_contents[14'h2f83] = 8'hdd;
s_mem_contents[14'h2f84] = 8'h62;
s_mem_contents[14'h2f85] = 8'h02;
s_mem_contents[14'h2f86] = 8'hd0;
s_mem_contents[14'h2f87] = 8'hfe;
s_mem_contents[14'h2f88] = 8'h68;
s_mem_contents[14'h2f89] = 8'h49;
s_mem_contents[14'h2f8a] = 8'h7d;
s_mem_contents[14'h2f8b] = 8'hdd;
s_mem_contents[14'h2f8c] = 8'h66;
s_mem_contents[14'h2f8d] = 8'h02;
s_mem_contents[14'h2f8e] = 8'hd0;
s_mem_contents[14'h2f8f] = 8'hfe;
s_mem_contents[14'h2f90] = 8'hca;
s_mem_contents[14'h2f91] = 8'h10;
s_mem_contents[14'h2f92] = 8'h02;
s_mem_contents[14'h2f93] = 8'ha2;
s_mem_contents[14'h2f94] = 8'h03;
s_mem_contents[14'h2f95] = 8'ha9;
s_mem_contents[14'h2f96] = 8'h00;
s_mem_contents[14'h2f97] = 8'h48;
s_mem_contents[14'h2f98] = 8'hbd;
s_mem_contents[14'h2f99] = 8'h5e;
s_mem_contents[14'h2f9a] = 8'h02;
s_mem_contents[14'h2f9b] = 8'h28;
s_mem_contents[14'h2f9c] = 8'h55;
s_mem_contents[14'h2f9d] = 8'h16;
s_mem_contents[14'h2f9e] = 8'h08;
s_mem_contents[14'h2f9f] = 8'hdd;
s_mem_contents[14'h2fa0] = 8'h62;
s_mem_contents[14'h2fa1] = 8'h02;
s_mem_contents[14'h2fa2] = 8'hd0;
s_mem_contents[14'h2fa3] = 8'hfe;
s_mem_contents[14'h2fa4] = 8'h68;
s_mem_contents[14'h2fa5] = 8'h49;
s_mem_contents[14'h2fa6] = 8'h30;
s_mem_contents[14'h2fa7] = 8'hdd;
s_mem_contents[14'h2fa8] = 8'h66;
s_mem_contents[14'h2fa9] = 8'h02;
s_mem_contents[14'h2faa] = 8'hd0;
s_mem_contents[14'h2fab] = 8'hfe;
s_mem_contents[14'h2fac] = 8'hca;
s_mem_contents[14'h2fad] = 8'h10;
s_mem_contents[14'h2fae] = 8'he6;
s_mem_contents[14'h2faf] = 8'ha2;
s_mem_contents[14'h2fb0] = 8'h03;
s_mem_contents[14'h2fb1] = 8'ha9;
s_mem_contents[14'h2fb2] = 8'hff;
s_mem_contents[14'h2fb3] = 8'h48;
s_mem_contents[14'h2fb4] = 8'hbd;
s_mem_contents[14'h2fb5] = 8'h5e;
s_mem_contents[14'h2fb6] = 8'h02;
s_mem_contents[14'h2fb7] = 8'h28;
s_mem_contents[14'h2fb8] = 8'h55;
s_mem_contents[14'h2fb9] = 8'h16;
s_mem_contents[14'h2fba] = 8'h08;
s_mem_contents[14'h2fbb] = 8'hdd;
s_mem_contents[14'h2fbc] = 8'h62;
s_mem_contents[14'h2fbd] = 8'h02;
s_mem_contents[14'h2fbe] = 8'hd0;
s_mem_contents[14'h2fbf] = 8'hfe;
s_mem_contents[14'h2fc0] = 8'h68;
s_mem_contents[14'h2fc1] = 8'h49;
s_mem_contents[14'h2fc2] = 8'h7d;
s_mem_contents[14'h2fc3] = 8'hdd;
s_mem_contents[14'h2fc4] = 8'h66;
s_mem_contents[14'h2fc5] = 8'h02;
s_mem_contents[14'h2fc6] = 8'hd0;
s_mem_contents[14'h2fc7] = 8'hfe;
s_mem_contents[14'h2fc8] = 8'hca;
s_mem_contents[14'h2fc9] = 8'h10;
s_mem_contents[14'h2fca] = 8'he6;
s_mem_contents[14'h2fcb] = 8'ha2;
s_mem_contents[14'h2fcc] = 8'h03;
s_mem_contents[14'h2fcd] = 8'ha9;
s_mem_contents[14'h2fce] = 8'h00;
s_mem_contents[14'h2fcf] = 8'h48;
s_mem_contents[14'h2fd0] = 8'hbd;
s_mem_contents[14'h2fd1] = 8'h5e;
s_mem_contents[14'h2fd2] = 8'h02;
s_mem_contents[14'h2fd3] = 8'h28;
s_mem_contents[14'h2fd4] = 8'h5d;
s_mem_contents[14'h2fd5] = 8'h52;
s_mem_contents[14'h2fd6] = 8'h02;
s_mem_contents[14'h2fd7] = 8'h08;
s_mem_contents[14'h2fd8] = 8'hdd;
s_mem_contents[14'h2fd9] = 8'h62;
s_mem_contents[14'h2fda] = 8'h02;
s_mem_contents[14'h2fdb] = 8'hd0;
s_mem_contents[14'h2fdc] = 8'hfe;
s_mem_contents[14'h2fdd] = 8'h68;
s_mem_contents[14'h2fde] = 8'h49;
s_mem_contents[14'h2fdf] = 8'h30;
s_mem_contents[14'h2fe0] = 8'hdd;
s_mem_contents[14'h2fe1] = 8'h66;
s_mem_contents[14'h2fe2] = 8'h02;
s_mem_contents[14'h2fe3] = 8'hd0;
s_mem_contents[14'h2fe4] = 8'hfe;
s_mem_contents[14'h2fe5] = 8'hca;
s_mem_contents[14'h2fe6] = 8'h10;
s_mem_contents[14'h2fe7] = 8'he5;
s_mem_contents[14'h2fe8] = 8'ha2;
s_mem_contents[14'h2fe9] = 8'h03;
s_mem_contents[14'h2fea] = 8'ha9;
s_mem_contents[14'h2feb] = 8'hff;
s_mem_contents[14'h2fec] = 8'h48;
s_mem_contents[14'h2fed] = 8'hbd;
s_mem_contents[14'h2fee] = 8'h5e;
s_mem_contents[14'h2fef] = 8'h02;
s_mem_contents[14'h2ff0] = 8'h28;
s_mem_contents[14'h2ff1] = 8'h5d;
s_mem_contents[14'h2ff2] = 8'h52;
s_mem_contents[14'h2ff3] = 8'h02;
s_mem_contents[14'h2ff4] = 8'h08;
s_mem_contents[14'h2ff5] = 8'hdd;
s_mem_contents[14'h2ff6] = 8'h62;
s_mem_contents[14'h2ff7] = 8'h02;
s_mem_contents[14'h2ff8] = 8'hd0;
s_mem_contents[14'h2ff9] = 8'hfe;
s_mem_contents[14'h2ffa] = 8'h68;
s_mem_contents[14'h2ffb] = 8'h49;
s_mem_contents[14'h2ffc] = 8'h7d;
s_mem_contents[14'h2ffd] = 8'hdd;
s_mem_contents[14'h2ffe] = 8'h66;
s_mem_contents[14'h2fff] = 8'h02;
s_mem_contents[14'h3000] = 8'hd0;
s_mem_contents[14'h3001] = 8'hfe;
s_mem_contents[14'h3002] = 8'hca;
s_mem_contents[14'h3003] = 8'h10;
s_mem_contents[14'h3004] = 8'he5;
s_mem_contents[14'h3005] = 8'ha0;
s_mem_contents[14'h3006] = 8'h03;
s_mem_contents[14'h3007] = 8'ha9;
s_mem_contents[14'h3008] = 8'h00;
s_mem_contents[14'h3009] = 8'h48;
s_mem_contents[14'h300a] = 8'hb9;
s_mem_contents[14'h300b] = 8'h5e;
s_mem_contents[14'h300c] = 8'h02;
s_mem_contents[14'h300d] = 8'h28;
s_mem_contents[14'h300e] = 8'h59;
s_mem_contents[14'h300f] = 8'h52;
s_mem_contents[14'h3010] = 8'h02;
s_mem_contents[14'h3011] = 8'h08;
s_mem_contents[14'h3012] = 8'hd9;
s_mem_contents[14'h3013] = 8'h62;
s_mem_contents[14'h3014] = 8'h02;
s_mem_contents[14'h3015] = 8'hd0;
s_mem_contents[14'h3016] = 8'hfe;
s_mem_contents[14'h3017] = 8'h68;
s_mem_contents[14'h3018] = 8'h49;
s_mem_contents[14'h3019] = 8'h30;
s_mem_contents[14'h301a] = 8'hd9;
s_mem_contents[14'h301b] = 8'h66;
s_mem_contents[14'h301c] = 8'h02;
s_mem_contents[14'h301d] = 8'hd0;
s_mem_contents[14'h301e] = 8'hfe;
s_mem_contents[14'h301f] = 8'h88;
s_mem_contents[14'h3020] = 8'h10;
s_mem_contents[14'h3021] = 8'he5;
s_mem_contents[14'h3022] = 8'ha0;
s_mem_contents[14'h3023] = 8'h03;
s_mem_contents[14'h3024] = 8'ha9;
s_mem_contents[14'h3025] = 8'hff;
s_mem_contents[14'h3026] = 8'h48;
s_mem_contents[14'h3027] = 8'hb9;
s_mem_contents[14'h3028] = 8'h5e;
s_mem_contents[14'h3029] = 8'h02;
s_mem_contents[14'h302a] = 8'h28;
s_mem_contents[14'h302b] = 8'h59;
s_mem_contents[14'h302c] = 8'h52;
s_mem_contents[14'h302d] = 8'h02;
s_mem_contents[14'h302e] = 8'h08;
s_mem_contents[14'h302f] = 8'hd9;
s_mem_contents[14'h3030] = 8'h62;
s_mem_contents[14'h3031] = 8'h02;
s_mem_contents[14'h3032] = 8'hd0;
s_mem_contents[14'h3033] = 8'hfe;
s_mem_contents[14'h3034] = 8'h68;
s_mem_contents[14'h3035] = 8'h49;
s_mem_contents[14'h3036] = 8'h7d;
s_mem_contents[14'h3037] = 8'hd9;
s_mem_contents[14'h3038] = 8'h66;
s_mem_contents[14'h3039] = 8'h02;
s_mem_contents[14'h303a] = 8'hd0;
s_mem_contents[14'h303b] = 8'hfe;
s_mem_contents[14'h303c] = 8'h88;
s_mem_contents[14'h303d] = 8'h10;
s_mem_contents[14'h303e] = 8'he5;
s_mem_contents[14'h303f] = 8'ha2;
s_mem_contents[14'h3040] = 8'h06;
s_mem_contents[14'h3041] = 8'ha0;
s_mem_contents[14'h3042] = 8'h03;
s_mem_contents[14'h3043] = 8'ha9;
s_mem_contents[14'h3044] = 8'h00;
s_mem_contents[14'h3045] = 8'h48;
s_mem_contents[14'h3046] = 8'hb9;
s_mem_contents[14'h3047] = 8'h5e;
s_mem_contents[14'h3048] = 8'h02;
s_mem_contents[14'h3049] = 8'h28;
s_mem_contents[14'h304a] = 8'h41;
s_mem_contents[14'h304b] = 8'h38;
s_mem_contents[14'h304c] = 8'h08;
s_mem_contents[14'h304d] = 8'hd9;
s_mem_contents[14'h304e] = 8'h62;
s_mem_contents[14'h304f] = 8'h02;
s_mem_contents[14'h3050] = 8'hd0;
s_mem_contents[14'h3051] = 8'hfe;
s_mem_contents[14'h3052] = 8'h68;
s_mem_contents[14'h3053] = 8'h49;
s_mem_contents[14'h3054] = 8'h30;
s_mem_contents[14'h3055] = 8'hd9;
s_mem_contents[14'h3056] = 8'h66;
s_mem_contents[14'h3057] = 8'h02;
s_mem_contents[14'h3058] = 8'hd0;
s_mem_contents[14'h3059] = 8'hfe;
s_mem_contents[14'h305a] = 8'hca;
s_mem_contents[14'h305b] = 8'hca;
s_mem_contents[14'h305c] = 8'h88;
s_mem_contents[14'h305d] = 8'h10;
s_mem_contents[14'h305e] = 8'he4;
s_mem_contents[14'h305f] = 8'ha2;
s_mem_contents[14'h3060] = 8'h06;
s_mem_contents[14'h3061] = 8'ha0;
s_mem_contents[14'h3062] = 8'h03;
s_mem_contents[14'h3063] = 8'ha9;
s_mem_contents[14'h3064] = 8'hff;
s_mem_contents[14'h3065] = 8'h48;
s_mem_contents[14'h3066] = 8'hb9;
s_mem_contents[14'h3067] = 8'h5e;
s_mem_contents[14'h3068] = 8'h02;
s_mem_contents[14'h3069] = 8'h28;
s_mem_contents[14'h306a] = 8'h41;
s_mem_contents[14'h306b] = 8'h38;
s_mem_contents[14'h306c] = 8'h08;
s_mem_contents[14'h306d] = 8'hd9;
s_mem_contents[14'h306e] = 8'h62;
s_mem_contents[14'h306f] = 8'h02;
s_mem_contents[14'h3070] = 8'hd0;
s_mem_contents[14'h3071] = 8'hfe;
s_mem_contents[14'h3072] = 8'h68;
s_mem_contents[14'h3073] = 8'h49;
s_mem_contents[14'h3074] = 8'h7d;
s_mem_contents[14'h3075] = 8'hd9;
s_mem_contents[14'h3076] = 8'h66;
s_mem_contents[14'h3077] = 8'h02;
s_mem_contents[14'h3078] = 8'hd0;
s_mem_contents[14'h3079] = 8'hfe;
s_mem_contents[14'h307a] = 8'hca;
s_mem_contents[14'h307b] = 8'hca;
s_mem_contents[14'h307c] = 8'h88;
s_mem_contents[14'h307d] = 8'h10;
s_mem_contents[14'h307e] = 8'he4;
s_mem_contents[14'h307f] = 8'ha0;
s_mem_contents[14'h3080] = 8'h03;
s_mem_contents[14'h3081] = 8'ha9;
s_mem_contents[14'h3082] = 8'h00;
s_mem_contents[14'h3083] = 8'h48;
s_mem_contents[14'h3084] = 8'hb9;
s_mem_contents[14'h3085] = 8'h5e;
s_mem_contents[14'h3086] = 8'h02;
s_mem_contents[14'h3087] = 8'h28;
s_mem_contents[14'h3088] = 8'h51;
s_mem_contents[14'h3089] = 8'h38;
s_mem_contents[14'h308a] = 8'h08;
s_mem_contents[14'h308b] = 8'hd9;
s_mem_contents[14'h308c] = 8'h62;
s_mem_contents[14'h308d] = 8'h02;
s_mem_contents[14'h308e] = 8'hd0;
s_mem_contents[14'h308f] = 8'hfe;
s_mem_contents[14'h3090] = 8'h68;
s_mem_contents[14'h3091] = 8'h49;
s_mem_contents[14'h3092] = 8'h30;
s_mem_contents[14'h3093] = 8'hd9;
s_mem_contents[14'h3094] = 8'h66;
s_mem_contents[14'h3095] = 8'h02;
s_mem_contents[14'h3096] = 8'hd0;
s_mem_contents[14'h3097] = 8'hfe;
s_mem_contents[14'h3098] = 8'h88;
s_mem_contents[14'h3099] = 8'h10;
s_mem_contents[14'h309a] = 8'he6;
s_mem_contents[14'h309b] = 8'ha0;
s_mem_contents[14'h309c] = 8'h03;
s_mem_contents[14'h309d] = 8'ha9;
s_mem_contents[14'h309e] = 8'hff;
s_mem_contents[14'h309f] = 8'h48;
s_mem_contents[14'h30a0] = 8'hb9;
s_mem_contents[14'h30a1] = 8'h5e;
s_mem_contents[14'h30a2] = 8'h02;
s_mem_contents[14'h30a3] = 8'h28;
s_mem_contents[14'h30a4] = 8'h51;
s_mem_contents[14'h30a5] = 8'h38;
s_mem_contents[14'h30a6] = 8'h08;
s_mem_contents[14'h30a7] = 8'hd9;
s_mem_contents[14'h30a8] = 8'h62;
s_mem_contents[14'h30a9] = 8'h02;
s_mem_contents[14'h30aa] = 8'hd0;
s_mem_contents[14'h30ab] = 8'hfe;
s_mem_contents[14'h30ac] = 8'h68;
s_mem_contents[14'h30ad] = 8'h49;
s_mem_contents[14'h30ae] = 8'h7d;
s_mem_contents[14'h30af] = 8'hd9;
s_mem_contents[14'h30b0] = 8'h66;
s_mem_contents[14'h30b1] = 8'h02;
s_mem_contents[14'h30b2] = 8'hd0;
s_mem_contents[14'h30b3] = 8'hfe;
s_mem_contents[14'h30b4] = 8'h88;
s_mem_contents[14'h30b5] = 8'h10;
s_mem_contents[14'h30b6] = 8'he6;
s_mem_contents[14'h30b7] = 8'had;
s_mem_contents[14'h30b8] = 8'h00;
s_mem_contents[14'h30b9] = 8'h02;
s_mem_contents[14'h30ba] = 8'hc9;
s_mem_contents[14'h30bb] = 8'h27;
s_mem_contents[14'h30bc] = 8'hd0;
s_mem_contents[14'h30bd] = 8'hfe;
s_mem_contents[14'h30be] = 8'ha9;
s_mem_contents[14'h30bf] = 8'h28;
s_mem_contents[14'h30c0] = 8'h8d;
s_mem_contents[14'h30c1] = 8'h00;
s_mem_contents[14'h30c2] = 8'h02;
s_mem_contents[14'h30c3] = 8'ha2;
s_mem_contents[14'h30c4] = 8'h03;
s_mem_contents[14'h30c5] = 8'hb5;
s_mem_contents[14'h30c6] = 8'h0e;
s_mem_contents[14'h30c7] = 8'h8d;
s_mem_contents[14'h30c8] = 8'h0f;
s_mem_contents[14'h30c9] = 8'h02;
s_mem_contents[14'h30ca] = 8'ha9;
s_mem_contents[14'h30cb] = 8'h00;
s_mem_contents[14'h30cc] = 8'h48;
s_mem_contents[14'h30cd] = 8'hbd;
s_mem_contents[14'h30ce] = 8'h56;
s_mem_contents[14'h30cf] = 8'h02;
s_mem_contents[14'h30d0] = 8'h28;
s_mem_contents[14'h30d1] = 8'h20;
s_mem_contents[14'h30d2] = 8'h0e;
s_mem_contents[14'h30d3] = 8'h02;
s_mem_contents[14'h30d4] = 8'h08;
s_mem_contents[14'h30d5] = 8'hdd;
s_mem_contents[14'h30d6] = 8'h62;
s_mem_contents[14'h30d7] = 8'h02;
s_mem_contents[14'h30d8] = 8'hd0;
s_mem_contents[14'h30d9] = 8'hfe;
s_mem_contents[14'h30da] = 8'h68;
s_mem_contents[14'h30db] = 8'h49;
s_mem_contents[14'h30dc] = 8'h30;
s_mem_contents[14'h30dd] = 8'hdd;
s_mem_contents[14'h30de] = 8'h66;
s_mem_contents[14'h30df] = 8'h02;
s_mem_contents[14'h30e0] = 8'hd0;
s_mem_contents[14'h30e1] = 8'hfe;
s_mem_contents[14'h30e2] = 8'hca;
s_mem_contents[14'h30e3] = 8'h10;
s_mem_contents[14'h30e4] = 8'he0;
s_mem_contents[14'h30e5] = 8'ha2;
s_mem_contents[14'h30e6] = 8'h03;
s_mem_contents[14'h30e7] = 8'hb5;
s_mem_contents[14'h30e8] = 8'h0e;
s_mem_contents[14'h30e9] = 8'h8d;
s_mem_contents[14'h30ea] = 8'h0f;
s_mem_contents[14'h30eb] = 8'h02;
s_mem_contents[14'h30ec] = 8'ha9;
s_mem_contents[14'h30ed] = 8'hff;
s_mem_contents[14'h30ee] = 8'h48;
s_mem_contents[14'h30ef] = 8'hbd;
s_mem_contents[14'h30f0] = 8'h56;
s_mem_contents[14'h30f1] = 8'h02;
s_mem_contents[14'h30f2] = 8'h28;
s_mem_contents[14'h30f3] = 8'h20;
s_mem_contents[14'h30f4] = 8'h0e;
s_mem_contents[14'h30f5] = 8'h02;
s_mem_contents[14'h30f6] = 8'h08;
s_mem_contents[14'h30f7] = 8'hdd;
s_mem_contents[14'h30f8] = 8'h62;
s_mem_contents[14'h30f9] = 8'h02;
s_mem_contents[14'h30fa] = 8'hd0;
s_mem_contents[14'h30fb] = 8'hfe;
s_mem_contents[14'h30fc] = 8'h68;
s_mem_contents[14'h30fd] = 8'h49;
s_mem_contents[14'h30fe] = 8'h7d;
s_mem_contents[14'h30ff] = 8'hdd;
s_mem_contents[14'h3100] = 8'h66;
s_mem_contents[14'h3101] = 8'h02;
s_mem_contents[14'h3102] = 8'hd0;
s_mem_contents[14'h3103] = 8'hfe;
s_mem_contents[14'h3104] = 8'hca;
s_mem_contents[14'h3105] = 8'h10;
s_mem_contents[14'h3106] = 8'he0;
s_mem_contents[14'h3107] = 8'ha2;
s_mem_contents[14'h3108] = 8'h03;
s_mem_contents[14'h3109] = 8'hb5;
s_mem_contents[14'h310a] = 8'h0e;
s_mem_contents[14'h310b] = 8'h85;
s_mem_contents[14'h310c] = 8'h02;
s_mem_contents[14'h310d] = 8'ha9;
s_mem_contents[14'h310e] = 8'h00;
s_mem_contents[14'h310f] = 8'h48;
s_mem_contents[14'h3110] = 8'hbd;
s_mem_contents[14'h3111] = 8'h56;
s_mem_contents[14'h3112] = 8'h02;
s_mem_contents[14'h3113] = 8'h28;
s_mem_contents[14'h3114] = 8'h05;
s_mem_contents[14'h3115] = 8'h02;
s_mem_contents[14'h3116] = 8'h08;
s_mem_contents[14'h3117] = 8'hdd;
s_mem_contents[14'h3118] = 8'h62;
s_mem_contents[14'h3119] = 8'h02;
s_mem_contents[14'h311a] = 8'hd0;
s_mem_contents[14'h311b] = 8'hfe;
s_mem_contents[14'h311c] = 8'h68;
s_mem_contents[14'h311d] = 8'h49;
s_mem_contents[14'h311e] = 8'h30;
s_mem_contents[14'h311f] = 8'hdd;
s_mem_contents[14'h3120] = 8'h66;
s_mem_contents[14'h3121] = 8'h02;
s_mem_contents[14'h3122] = 8'hd0;
s_mem_contents[14'h3123] = 8'hfe;
s_mem_contents[14'h3124] = 8'hca;
s_mem_contents[14'h3125] = 8'h10;
s_mem_contents[14'h3126] = 8'he2;
s_mem_contents[14'h3127] = 8'ha2;
s_mem_contents[14'h3128] = 8'h03;
s_mem_contents[14'h3129] = 8'hb5;
s_mem_contents[14'h312a] = 8'h0e;
s_mem_contents[14'h312b] = 8'h85;
s_mem_contents[14'h312c] = 8'h02;
s_mem_contents[14'h312d] = 8'ha9;
s_mem_contents[14'h312e] = 8'hff;
s_mem_contents[14'h312f] = 8'h48;
s_mem_contents[14'h3130] = 8'hbd;
s_mem_contents[14'h3131] = 8'h56;
s_mem_contents[14'h3132] = 8'h02;
s_mem_contents[14'h3133] = 8'h28;
s_mem_contents[14'h3134] = 8'h05;
s_mem_contents[14'h3135] = 8'h02;
s_mem_contents[14'h3136] = 8'h08;
s_mem_contents[14'h3137] = 8'hdd;
s_mem_contents[14'h3138] = 8'h62;
s_mem_contents[14'h3139] = 8'h02;
s_mem_contents[14'h313a] = 8'hd0;
s_mem_contents[14'h313b] = 8'hfe;
s_mem_contents[14'h313c] = 8'h68;
s_mem_contents[14'h313d] = 8'h49;
s_mem_contents[14'h313e] = 8'h7d;
s_mem_contents[14'h313f] = 8'hdd;
s_mem_contents[14'h3140] = 8'h66;
s_mem_contents[14'h3141] = 8'h02;
s_mem_contents[14'h3142] = 8'hd0;
s_mem_contents[14'h3143] = 8'hfe;
s_mem_contents[14'h3144] = 8'hca;
s_mem_contents[14'h3145] = 8'h10;
s_mem_contents[14'h3146] = 8'he2;
s_mem_contents[14'h3147] = 8'ha2;
s_mem_contents[14'h3148] = 8'h03;
s_mem_contents[14'h3149] = 8'hb5;
s_mem_contents[14'h314a] = 8'h0e;
s_mem_contents[14'h314b] = 8'h8d;
s_mem_contents[14'h314c] = 8'h03;
s_mem_contents[14'h314d] = 8'h02;
s_mem_contents[14'h314e] = 8'ha9;
s_mem_contents[14'h314f] = 8'h00;
s_mem_contents[14'h3150] = 8'h48;
s_mem_contents[14'h3151] = 8'hbd;
s_mem_contents[14'h3152] = 8'h56;
s_mem_contents[14'h3153] = 8'h02;
s_mem_contents[14'h3154] = 8'h28;
s_mem_contents[14'h3155] = 8'h0d;
s_mem_contents[14'h3156] = 8'h03;
s_mem_contents[14'h3157] = 8'h02;
s_mem_contents[14'h3158] = 8'h08;
s_mem_contents[14'h3159] = 8'hdd;
s_mem_contents[14'h315a] = 8'h62;
s_mem_contents[14'h315b] = 8'h02;
s_mem_contents[14'h315c] = 8'hd0;
s_mem_contents[14'h315d] = 8'hfe;
s_mem_contents[14'h315e] = 8'h68;
s_mem_contents[14'h315f] = 8'h49;
s_mem_contents[14'h3160] = 8'h30;
s_mem_contents[14'h3161] = 8'hdd;
s_mem_contents[14'h3162] = 8'h66;
s_mem_contents[14'h3163] = 8'h02;
s_mem_contents[14'h3164] = 8'hd0;
s_mem_contents[14'h3165] = 8'hfe;
s_mem_contents[14'h3166] = 8'hca;
s_mem_contents[14'h3167] = 8'h10;
s_mem_contents[14'h3168] = 8'he0;
s_mem_contents[14'h3169] = 8'ha2;
s_mem_contents[14'h316a] = 8'h03;
s_mem_contents[14'h316b] = 8'hb5;
s_mem_contents[14'h316c] = 8'h0e;
s_mem_contents[14'h316d] = 8'h8d;
s_mem_contents[14'h316e] = 8'h03;
s_mem_contents[14'h316f] = 8'h02;
s_mem_contents[14'h3170] = 8'ha9;
s_mem_contents[14'h3171] = 8'hff;
s_mem_contents[14'h3172] = 8'h48;
s_mem_contents[14'h3173] = 8'hbd;
s_mem_contents[14'h3174] = 8'h56;
s_mem_contents[14'h3175] = 8'h02;
s_mem_contents[14'h3176] = 8'h28;
s_mem_contents[14'h3177] = 8'h0d;
s_mem_contents[14'h3178] = 8'h03;
s_mem_contents[14'h3179] = 8'h02;
s_mem_contents[14'h317a] = 8'h08;
s_mem_contents[14'h317b] = 8'hdd;
s_mem_contents[14'h317c] = 8'h62;
s_mem_contents[14'h317d] = 8'h02;
s_mem_contents[14'h317e] = 8'hd0;
s_mem_contents[14'h317f] = 8'hfe;
s_mem_contents[14'h3180] = 8'h68;
s_mem_contents[14'h3181] = 8'h49;
s_mem_contents[14'h3182] = 8'h7d;
s_mem_contents[14'h3183] = 8'hdd;
s_mem_contents[14'h3184] = 8'h66;
s_mem_contents[14'h3185] = 8'h02;
s_mem_contents[14'h3186] = 8'hd0;
s_mem_contents[14'h3187] = 8'hfe;
s_mem_contents[14'h3188] = 8'hca;
s_mem_contents[14'h3189] = 8'h10;
s_mem_contents[14'h318a] = 8'h02;
s_mem_contents[14'h318b] = 8'ha2;
s_mem_contents[14'h318c] = 8'h03;
s_mem_contents[14'h318d] = 8'ha9;
s_mem_contents[14'h318e] = 8'h00;
s_mem_contents[14'h318f] = 8'h48;
s_mem_contents[14'h3190] = 8'hbd;
s_mem_contents[14'h3191] = 8'h56;
s_mem_contents[14'h3192] = 8'h02;
s_mem_contents[14'h3193] = 8'h28;
s_mem_contents[14'h3194] = 8'h15;
s_mem_contents[14'h3195] = 8'h0e;
s_mem_contents[14'h3196] = 8'h08;
s_mem_contents[14'h3197] = 8'hdd;
s_mem_contents[14'h3198] = 8'h62;
s_mem_contents[14'h3199] = 8'h02;
s_mem_contents[14'h319a] = 8'hd0;
s_mem_contents[14'h319b] = 8'hfe;
s_mem_contents[14'h319c] = 8'h68;
s_mem_contents[14'h319d] = 8'h49;
s_mem_contents[14'h319e] = 8'h30;
s_mem_contents[14'h319f] = 8'hdd;
s_mem_contents[14'h31a0] = 8'h66;
s_mem_contents[14'h31a1] = 8'h02;
s_mem_contents[14'h31a2] = 8'hd0;
s_mem_contents[14'h31a3] = 8'hfe;
s_mem_contents[14'h31a4] = 8'hca;
s_mem_contents[14'h31a5] = 8'h10;
s_mem_contents[14'h31a6] = 8'he6;
s_mem_contents[14'h31a7] = 8'ha2;
s_mem_contents[14'h31a8] = 8'h03;
s_mem_contents[14'h31a9] = 8'ha9;
s_mem_contents[14'h31aa] = 8'hff;
s_mem_contents[14'h31ab] = 8'h48;
s_mem_contents[14'h31ac] = 8'hbd;
s_mem_contents[14'h31ad] = 8'h56;
s_mem_contents[14'h31ae] = 8'h02;
s_mem_contents[14'h31af] = 8'h28;
s_mem_contents[14'h31b0] = 8'h15;
s_mem_contents[14'h31b1] = 8'h0e;
s_mem_contents[14'h31b2] = 8'h08;
s_mem_contents[14'h31b3] = 8'hdd;
s_mem_contents[14'h31b4] = 8'h62;
s_mem_contents[14'h31b5] = 8'h02;
s_mem_contents[14'h31b6] = 8'hd0;
s_mem_contents[14'h31b7] = 8'hfe;
s_mem_contents[14'h31b8] = 8'h68;
s_mem_contents[14'h31b9] = 8'h49;
s_mem_contents[14'h31ba] = 8'h7d;
s_mem_contents[14'h31bb] = 8'hdd;
s_mem_contents[14'h31bc] = 8'h66;
s_mem_contents[14'h31bd] = 8'h02;
s_mem_contents[14'h31be] = 8'hd0;
s_mem_contents[14'h31bf] = 8'hfe;
s_mem_contents[14'h31c0] = 8'hca;
s_mem_contents[14'h31c1] = 8'h10;
s_mem_contents[14'h31c2] = 8'he6;
s_mem_contents[14'h31c3] = 8'ha2;
s_mem_contents[14'h31c4] = 8'h03;
s_mem_contents[14'h31c5] = 8'ha9;
s_mem_contents[14'h31c6] = 8'h00;
s_mem_contents[14'h31c7] = 8'h48;
s_mem_contents[14'h31c8] = 8'hbd;
s_mem_contents[14'h31c9] = 8'h56;
s_mem_contents[14'h31ca] = 8'h02;
s_mem_contents[14'h31cb] = 8'h28;
s_mem_contents[14'h31cc] = 8'h1d;
s_mem_contents[14'h31cd] = 8'h4a;
s_mem_contents[14'h31ce] = 8'h02;
s_mem_contents[14'h31cf] = 8'h08;
s_mem_contents[14'h31d0] = 8'hdd;
s_mem_contents[14'h31d1] = 8'h62;
s_mem_contents[14'h31d2] = 8'h02;
s_mem_contents[14'h31d3] = 8'hd0;
s_mem_contents[14'h31d4] = 8'hfe;
s_mem_contents[14'h31d5] = 8'h68;
s_mem_contents[14'h31d6] = 8'h49;
s_mem_contents[14'h31d7] = 8'h30;
s_mem_contents[14'h31d8] = 8'hdd;
s_mem_contents[14'h31d9] = 8'h66;
s_mem_contents[14'h31da] = 8'h02;
s_mem_contents[14'h31db] = 8'hd0;
s_mem_contents[14'h31dc] = 8'hfe;
s_mem_contents[14'h31dd] = 8'hca;
s_mem_contents[14'h31de] = 8'h10;
s_mem_contents[14'h31df] = 8'he5;
s_mem_contents[14'h31e0] = 8'ha2;
s_mem_contents[14'h31e1] = 8'h03;
s_mem_contents[14'h31e2] = 8'ha9;
s_mem_contents[14'h31e3] = 8'hff;
s_mem_contents[14'h31e4] = 8'h48;
s_mem_contents[14'h31e5] = 8'hbd;
s_mem_contents[14'h31e6] = 8'h56;
s_mem_contents[14'h31e7] = 8'h02;
s_mem_contents[14'h31e8] = 8'h28;
s_mem_contents[14'h31e9] = 8'h1d;
s_mem_contents[14'h31ea] = 8'h4a;
s_mem_contents[14'h31eb] = 8'h02;
s_mem_contents[14'h31ec] = 8'h08;
s_mem_contents[14'h31ed] = 8'hdd;
s_mem_contents[14'h31ee] = 8'h62;
s_mem_contents[14'h31ef] = 8'h02;
s_mem_contents[14'h31f0] = 8'hd0;
s_mem_contents[14'h31f1] = 8'hfe;
s_mem_contents[14'h31f2] = 8'h68;
s_mem_contents[14'h31f3] = 8'h49;
s_mem_contents[14'h31f4] = 8'h7d;
s_mem_contents[14'h31f5] = 8'hdd;
s_mem_contents[14'h31f6] = 8'h66;
s_mem_contents[14'h31f7] = 8'h02;
s_mem_contents[14'h31f8] = 8'hd0;
s_mem_contents[14'h31f9] = 8'hfe;
s_mem_contents[14'h31fa] = 8'hca;
s_mem_contents[14'h31fb] = 8'h10;
s_mem_contents[14'h31fc] = 8'he5;
s_mem_contents[14'h31fd] = 8'ha0;
s_mem_contents[14'h31fe] = 8'h03;
s_mem_contents[14'h31ff] = 8'ha9;
s_mem_contents[14'h3200] = 8'h00;
s_mem_contents[14'h3201] = 8'h48;
s_mem_contents[14'h3202] = 8'hb9;
s_mem_contents[14'h3203] = 8'h56;
s_mem_contents[14'h3204] = 8'h02;
s_mem_contents[14'h3205] = 8'h28;
s_mem_contents[14'h3206] = 8'h19;
s_mem_contents[14'h3207] = 8'h4a;
s_mem_contents[14'h3208] = 8'h02;
s_mem_contents[14'h3209] = 8'h08;
s_mem_contents[14'h320a] = 8'hd9;
s_mem_contents[14'h320b] = 8'h62;
s_mem_contents[14'h320c] = 8'h02;
s_mem_contents[14'h320d] = 8'hd0;
s_mem_contents[14'h320e] = 8'hfe;
s_mem_contents[14'h320f] = 8'h68;
s_mem_contents[14'h3210] = 8'h49;
s_mem_contents[14'h3211] = 8'h30;
s_mem_contents[14'h3212] = 8'hd9;
s_mem_contents[14'h3213] = 8'h66;
s_mem_contents[14'h3214] = 8'h02;
s_mem_contents[14'h3215] = 8'hd0;
s_mem_contents[14'h3216] = 8'hfe;
s_mem_contents[14'h3217] = 8'h88;
s_mem_contents[14'h3218] = 8'h10;
s_mem_contents[14'h3219] = 8'he5;
s_mem_contents[14'h321a] = 8'ha0;
s_mem_contents[14'h321b] = 8'h03;
s_mem_contents[14'h321c] = 8'ha9;
s_mem_contents[14'h321d] = 8'hff;
s_mem_contents[14'h321e] = 8'h48;
s_mem_contents[14'h321f] = 8'hb9;
s_mem_contents[14'h3220] = 8'h56;
s_mem_contents[14'h3221] = 8'h02;
s_mem_contents[14'h3222] = 8'h28;
s_mem_contents[14'h3223] = 8'h19;
s_mem_contents[14'h3224] = 8'h4a;
s_mem_contents[14'h3225] = 8'h02;
s_mem_contents[14'h3226] = 8'h08;
s_mem_contents[14'h3227] = 8'hd9;
s_mem_contents[14'h3228] = 8'h62;
s_mem_contents[14'h3229] = 8'h02;
s_mem_contents[14'h322a] = 8'hd0;
s_mem_contents[14'h322b] = 8'hfe;
s_mem_contents[14'h322c] = 8'h68;
s_mem_contents[14'h322d] = 8'h49;
s_mem_contents[14'h322e] = 8'h7d;
s_mem_contents[14'h322f] = 8'hd9;
s_mem_contents[14'h3230] = 8'h66;
s_mem_contents[14'h3231] = 8'h02;
s_mem_contents[14'h3232] = 8'hd0;
s_mem_contents[14'h3233] = 8'hfe;
s_mem_contents[14'h3234] = 8'h88;
s_mem_contents[14'h3235] = 8'h10;
s_mem_contents[14'h3236] = 8'he5;
s_mem_contents[14'h3237] = 8'ha2;
s_mem_contents[14'h3238] = 8'h06;
s_mem_contents[14'h3239] = 8'ha0;
s_mem_contents[14'h323a] = 8'h03;
s_mem_contents[14'h323b] = 8'ha9;
s_mem_contents[14'h323c] = 8'h00;
s_mem_contents[14'h323d] = 8'h48;
s_mem_contents[14'h323e] = 8'hb9;
s_mem_contents[14'h323f] = 8'h56;
s_mem_contents[14'h3240] = 8'h02;
s_mem_contents[14'h3241] = 8'h28;
s_mem_contents[14'h3242] = 8'h01;
s_mem_contents[14'h3243] = 8'h40;
s_mem_contents[14'h3244] = 8'h08;
s_mem_contents[14'h3245] = 8'hd9;
s_mem_contents[14'h3246] = 8'h62;
s_mem_contents[14'h3247] = 8'h02;
s_mem_contents[14'h3248] = 8'hd0;
s_mem_contents[14'h3249] = 8'hfe;
s_mem_contents[14'h324a] = 8'h68;
s_mem_contents[14'h324b] = 8'h49;
s_mem_contents[14'h324c] = 8'h30;
s_mem_contents[14'h324d] = 8'hd9;
s_mem_contents[14'h324e] = 8'h66;
s_mem_contents[14'h324f] = 8'h02;
s_mem_contents[14'h3250] = 8'hd0;
s_mem_contents[14'h3251] = 8'hfe;
s_mem_contents[14'h3252] = 8'hca;
s_mem_contents[14'h3253] = 8'hca;
s_mem_contents[14'h3254] = 8'h88;
s_mem_contents[14'h3255] = 8'h10;
s_mem_contents[14'h3256] = 8'he4;
s_mem_contents[14'h3257] = 8'ha2;
s_mem_contents[14'h3258] = 8'h06;
s_mem_contents[14'h3259] = 8'ha0;
s_mem_contents[14'h325a] = 8'h03;
s_mem_contents[14'h325b] = 8'ha9;
s_mem_contents[14'h325c] = 8'hff;
s_mem_contents[14'h325d] = 8'h48;
s_mem_contents[14'h325e] = 8'hb9;
s_mem_contents[14'h325f] = 8'h56;
s_mem_contents[14'h3260] = 8'h02;
s_mem_contents[14'h3261] = 8'h28;
s_mem_contents[14'h3262] = 8'h01;
s_mem_contents[14'h3263] = 8'h40;
s_mem_contents[14'h3264] = 8'h08;
s_mem_contents[14'h3265] = 8'hd9;
s_mem_contents[14'h3266] = 8'h62;
s_mem_contents[14'h3267] = 8'h02;
s_mem_contents[14'h3268] = 8'hd0;
s_mem_contents[14'h3269] = 8'hfe;
s_mem_contents[14'h326a] = 8'h68;
s_mem_contents[14'h326b] = 8'h49;
s_mem_contents[14'h326c] = 8'h7d;
s_mem_contents[14'h326d] = 8'hd9;
s_mem_contents[14'h326e] = 8'h66;
s_mem_contents[14'h326f] = 8'h02;
s_mem_contents[14'h3270] = 8'hd0;
s_mem_contents[14'h3271] = 8'hfe;
s_mem_contents[14'h3272] = 8'hca;
s_mem_contents[14'h3273] = 8'hca;
s_mem_contents[14'h3274] = 8'h88;
s_mem_contents[14'h3275] = 8'h10;
s_mem_contents[14'h3276] = 8'he4;
s_mem_contents[14'h3277] = 8'ha0;
s_mem_contents[14'h3278] = 8'h03;
s_mem_contents[14'h3279] = 8'ha9;
s_mem_contents[14'h327a] = 8'h00;
s_mem_contents[14'h327b] = 8'h48;
s_mem_contents[14'h327c] = 8'hb9;
s_mem_contents[14'h327d] = 8'h56;
s_mem_contents[14'h327e] = 8'h02;
s_mem_contents[14'h327f] = 8'h28;
s_mem_contents[14'h3280] = 8'h11;
s_mem_contents[14'h3281] = 8'h40;
s_mem_contents[14'h3282] = 8'h08;
s_mem_contents[14'h3283] = 8'hd9;
s_mem_contents[14'h3284] = 8'h62;
s_mem_contents[14'h3285] = 8'h02;
s_mem_contents[14'h3286] = 8'hd0;
s_mem_contents[14'h3287] = 8'hfe;
s_mem_contents[14'h3288] = 8'h68;
s_mem_contents[14'h3289] = 8'h49;
s_mem_contents[14'h328a] = 8'h30;
s_mem_contents[14'h328b] = 8'hd9;
s_mem_contents[14'h328c] = 8'h66;
s_mem_contents[14'h328d] = 8'h02;
s_mem_contents[14'h328e] = 8'hd0;
s_mem_contents[14'h328f] = 8'hfe;
s_mem_contents[14'h3290] = 8'h88;
s_mem_contents[14'h3291] = 8'h10;
s_mem_contents[14'h3292] = 8'he6;
s_mem_contents[14'h3293] = 8'ha0;
s_mem_contents[14'h3294] = 8'h03;
s_mem_contents[14'h3295] = 8'ha9;
s_mem_contents[14'h3296] = 8'hff;
s_mem_contents[14'h3297] = 8'h48;
s_mem_contents[14'h3298] = 8'hb9;
s_mem_contents[14'h3299] = 8'h56;
s_mem_contents[14'h329a] = 8'h02;
s_mem_contents[14'h329b] = 8'h28;
s_mem_contents[14'h329c] = 8'h11;
s_mem_contents[14'h329d] = 8'h40;
s_mem_contents[14'h329e] = 8'h08;
s_mem_contents[14'h329f] = 8'hd9;
s_mem_contents[14'h32a0] = 8'h62;
s_mem_contents[14'h32a1] = 8'h02;
s_mem_contents[14'h32a2] = 8'hd0;
s_mem_contents[14'h32a3] = 8'hfe;
s_mem_contents[14'h32a4] = 8'h68;
s_mem_contents[14'h32a5] = 8'h49;
s_mem_contents[14'h32a6] = 8'h7d;
s_mem_contents[14'h32a7] = 8'hd9;
s_mem_contents[14'h32a8] = 8'h66;
s_mem_contents[14'h32a9] = 8'h02;
s_mem_contents[14'h32aa] = 8'hd0;
s_mem_contents[14'h32ab] = 8'hfe;
s_mem_contents[14'h32ac] = 8'h88;
s_mem_contents[14'h32ad] = 8'h10;
s_mem_contents[14'h32ae] = 8'he6;
s_mem_contents[14'h32af] = 8'h58;
s_mem_contents[14'h32b0] = 8'had;
s_mem_contents[14'h32b1] = 8'h00;
s_mem_contents[14'h32b2] = 8'h02;
s_mem_contents[14'h32b3] = 8'hc9;
s_mem_contents[14'h32b4] = 8'h28;
s_mem_contents[14'h32b5] = 8'hd0;
s_mem_contents[14'h32b6] = 8'hfe;
s_mem_contents[14'h32b7] = 8'ha9;
s_mem_contents[14'h32b8] = 8'h29;
s_mem_contents[14'h32b9] = 8'h8d;
s_mem_contents[14'h32ba] = 8'h00;
s_mem_contents[14'h32bb] = 8'h02;
s_mem_contents[14'h32bc] = 8'hd8;
s_mem_contents[14'h32bd] = 8'ha2;
s_mem_contents[14'h32be] = 8'h04;
s_mem_contents[14'h32bf] = 8'ha0;
s_mem_contents[14'h32c0] = 8'hff;
s_mem_contents[14'h32c1] = 8'ha9;
s_mem_contents[14'h32c2] = 8'h00;
s_mem_contents[14'h32c3] = 8'h85;
s_mem_contents[14'h32c4] = 8'h02;
s_mem_contents[14'h32c5] = 8'h85;
s_mem_contents[14'h32c6] = 8'h03;
s_mem_contents[14'h32c7] = 8'h85;
s_mem_contents[14'h32c8] = 8'h04;
s_mem_contents[14'h32c9] = 8'h8d;
s_mem_contents[14'h32ca] = 8'h03;
s_mem_contents[14'h32cb] = 8'h02;
s_mem_contents[14'h32cc] = 8'h85;
s_mem_contents[14'h32cd] = 8'h05;
s_mem_contents[14'h32ce] = 8'h85;
s_mem_contents[14'h32cf] = 8'h06;
s_mem_contents[14'h32d0] = 8'ha9;
s_mem_contents[14'h32d1] = 8'hff;
s_mem_contents[14'h32d2] = 8'h85;
s_mem_contents[14'h32d3] = 8'h08;
s_mem_contents[14'h32d4] = 8'h8d;
s_mem_contents[14'h32d5] = 8'h04;
s_mem_contents[14'h32d6] = 8'h02;
s_mem_contents[14'h32d7] = 8'ha9;
s_mem_contents[14'h32d8] = 8'h02;
s_mem_contents[14'h32d9] = 8'h85;
s_mem_contents[14'h32da] = 8'h07;
s_mem_contents[14'h32db] = 8'h18;
s_mem_contents[14'h32dc] = 8'h20;
s_mem_contents[14'h32dd] = 8'h27;
s_mem_contents[14'h32de] = 8'h33;
s_mem_contents[14'h32df] = 8'he6;
s_mem_contents[14'h32e0] = 8'h02;
s_mem_contents[14'h32e1] = 8'he6;
s_mem_contents[14'h32e2] = 8'h05;
s_mem_contents[14'h32e3] = 8'h08;
s_mem_contents[14'h32e4] = 8'h08;
s_mem_contents[14'h32e5] = 8'h68;
s_mem_contents[14'h32e6] = 8'h29;
s_mem_contents[14'h32e7] = 8'h82;
s_mem_contents[14'h32e8] = 8'h28;
s_mem_contents[14'h32e9] = 8'hd0;
s_mem_contents[14'h32ea] = 8'h02;
s_mem_contents[14'h32eb] = 8'he6;
s_mem_contents[14'h32ec] = 8'h06;
s_mem_contents[14'h32ed] = 8'h05;
s_mem_contents[14'h32ee] = 8'h06;
s_mem_contents[14'h32ef] = 8'h85;
s_mem_contents[14'h32f0] = 8'h07;
s_mem_contents[14'h32f1] = 8'h38;
s_mem_contents[14'h32f2] = 8'h20;
s_mem_contents[14'h32f3] = 8'h27;
s_mem_contents[14'h32f4] = 8'h33;
s_mem_contents[14'h32f5] = 8'hc6;
s_mem_contents[14'h32f6] = 8'h02;
s_mem_contents[14'h32f7] = 8'he6;
s_mem_contents[14'h32f8] = 8'h03;
s_mem_contents[14'h32f9] = 8'hd0;
s_mem_contents[14'h32fa] = 8'he0;
s_mem_contents[14'h32fb] = 8'ha9;
s_mem_contents[14'h32fc] = 8'h00;
s_mem_contents[14'h32fd] = 8'h85;
s_mem_contents[14'h32fe] = 8'h06;
s_mem_contents[14'h32ff] = 8'hee;
s_mem_contents[14'h3300] = 8'h03;
s_mem_contents[14'h3301] = 8'h02;
s_mem_contents[14'h3302] = 8'he6;
s_mem_contents[14'h3303] = 8'h04;
s_mem_contents[14'h3304] = 8'h08;
s_mem_contents[14'h3305] = 8'h68;
s_mem_contents[14'h3306] = 8'h29;
s_mem_contents[14'h3307] = 8'h82;
s_mem_contents[14'h3308] = 8'h85;
s_mem_contents[14'h3309] = 8'h07;
s_mem_contents[14'h330a] = 8'hc6;
s_mem_contents[14'h330b] = 8'h08;
s_mem_contents[14'h330c] = 8'hce;
s_mem_contents[14'h330d] = 8'h04;
s_mem_contents[14'h330e] = 8'h02;
s_mem_contents[14'h330f] = 8'ha5;
s_mem_contents[14'h3310] = 8'h04;
s_mem_contents[14'h3311] = 8'h85;
s_mem_contents[14'h3312] = 8'h05;
s_mem_contents[14'h3313] = 8'hd0;
s_mem_contents[14'h3314] = 8'hc6;
s_mem_contents[14'h3315] = 8'had;
s_mem_contents[14'h3316] = 8'h00;
s_mem_contents[14'h3317] = 8'h02;
s_mem_contents[14'h3318] = 8'hc9;
s_mem_contents[14'h3319] = 8'h29;
s_mem_contents[14'h331a] = 8'hd0;
s_mem_contents[14'h331b] = 8'hfe;
s_mem_contents[14'h331c] = 8'ha9;
s_mem_contents[14'h331d] = 8'hf0;
s_mem_contents[14'h331e] = 8'h8d;
s_mem_contents[14'h331f] = 8'h00;
s_mem_contents[14'h3320] = 8'h02;
s_mem_contents[14'h3321] = 8'h4c;
s_mem_contents[14'h3322] = 8'h21;
s_mem_contents[14'h3323] = 8'h33;
s_mem_contents[14'h3324] = 8'h4c;
s_mem_contents[14'h3325] = 8'h00;
s_mem_contents[14'h3326] = 8'h04;
s_mem_contents[14'h3327] = 8'ha5;
s_mem_contents[14'h3328] = 8'h07;
s_mem_contents[14'h3329] = 8'h29;
s_mem_contents[14'h332a] = 8'h83;
s_mem_contents[14'h332b] = 8'h48;
s_mem_contents[14'h332c] = 8'ha5;
s_mem_contents[14'h332d] = 8'h03;
s_mem_contents[14'h332e] = 8'h45;
s_mem_contents[14'h332f] = 8'h04;
s_mem_contents[14'h3330] = 8'h30;
s_mem_contents[14'h3331] = 8'h0a;
s_mem_contents[14'h3332] = 8'ha5;
s_mem_contents[14'h3333] = 8'h03;
s_mem_contents[14'h3334] = 8'h45;
s_mem_contents[14'h3335] = 8'h05;
s_mem_contents[14'h3336] = 8'h10;
s_mem_contents[14'h3337] = 8'h04;
s_mem_contents[14'h3338] = 8'h68;
s_mem_contents[14'h3339] = 8'h09;
s_mem_contents[14'h333a] = 8'h40;
s_mem_contents[14'h333b] = 8'h48;
s_mem_contents[14'h333c] = 8'h68;
s_mem_contents[14'h333d] = 8'h85;
s_mem_contents[14'h333e] = 8'h07;
s_mem_contents[14'h333f] = 8'h08;
s_mem_contents[14'h3340] = 8'ha5;
s_mem_contents[14'h3341] = 8'h03;
s_mem_contents[14'h3342] = 8'h65;
s_mem_contents[14'h3343] = 8'h04;
s_mem_contents[14'h3344] = 8'h08;
s_mem_contents[14'h3345] = 8'hc5;
s_mem_contents[14'h3346] = 8'h05;
s_mem_contents[14'h3347] = 8'hd0;
s_mem_contents[14'h3348] = 8'hfe;
s_mem_contents[14'h3349] = 8'h68;
s_mem_contents[14'h334a] = 8'h29;
s_mem_contents[14'h334b] = 8'hc3;
s_mem_contents[14'h334c] = 8'hc5;
s_mem_contents[14'h334d] = 8'h07;
s_mem_contents[14'h334e] = 8'hd0;
s_mem_contents[14'h334f] = 8'hfe;
s_mem_contents[14'h3350] = 8'h28;
s_mem_contents[14'h3351] = 8'h08;
s_mem_contents[14'h3352] = 8'ha5;
s_mem_contents[14'h3353] = 8'h03;
s_mem_contents[14'h3354] = 8'he5;
s_mem_contents[14'h3355] = 8'h08;
s_mem_contents[14'h3356] = 8'h08;
s_mem_contents[14'h3357] = 8'hc5;
s_mem_contents[14'h3358] = 8'h05;
s_mem_contents[14'h3359] = 8'hd0;
s_mem_contents[14'h335a] = 8'hfe;
s_mem_contents[14'h335b] = 8'h68;
s_mem_contents[14'h335c] = 8'h29;
s_mem_contents[14'h335d] = 8'hc3;
s_mem_contents[14'h335e] = 8'hc5;
s_mem_contents[14'h335f] = 8'h07;
s_mem_contents[14'h3360] = 8'hd0;
s_mem_contents[14'h3361] = 8'hfe;
s_mem_contents[14'h3362] = 8'h28;
s_mem_contents[14'h3363] = 8'h08;
s_mem_contents[14'h3364] = 8'ha5;
s_mem_contents[14'h3365] = 8'h03;
s_mem_contents[14'h3366] = 8'h6d;
s_mem_contents[14'h3367] = 8'h03;
s_mem_contents[14'h3368] = 8'h02;
s_mem_contents[14'h3369] = 8'h08;
s_mem_contents[14'h336a] = 8'hc5;
s_mem_contents[14'h336b] = 8'h05;
s_mem_contents[14'h336c] = 8'hd0;
s_mem_contents[14'h336d] = 8'hfe;
s_mem_contents[14'h336e] = 8'h68;
s_mem_contents[14'h336f] = 8'h29;
s_mem_contents[14'h3370] = 8'hc3;
s_mem_contents[14'h3371] = 8'hc5;
s_mem_contents[14'h3372] = 8'h07;
s_mem_contents[14'h3373] = 8'hd0;
s_mem_contents[14'h3374] = 8'hfe;
s_mem_contents[14'h3375] = 8'h28;
s_mem_contents[14'h3376] = 8'h08;
s_mem_contents[14'h3377] = 8'ha5;
s_mem_contents[14'h3378] = 8'h03;
s_mem_contents[14'h3379] = 8'hed;
s_mem_contents[14'h337a] = 8'h04;
s_mem_contents[14'h337b] = 8'h02;
s_mem_contents[14'h337c] = 8'h08;
s_mem_contents[14'h337d] = 8'hc5;
s_mem_contents[14'h337e] = 8'h05;
s_mem_contents[14'h337f] = 8'hd0;
s_mem_contents[14'h3380] = 8'hfe;
s_mem_contents[14'h3381] = 8'h68;
s_mem_contents[14'h3382] = 8'h29;
s_mem_contents[14'h3383] = 8'hc3;
s_mem_contents[14'h3384] = 8'hc5;
s_mem_contents[14'h3385] = 8'h07;
s_mem_contents[14'h3386] = 8'hd0;
s_mem_contents[14'h3387] = 8'hfe;
s_mem_contents[14'h3388] = 8'h28;
s_mem_contents[14'h3389] = 8'h08;
s_mem_contents[14'h338a] = 8'ha5;
s_mem_contents[14'h338b] = 8'h04;
s_mem_contents[14'h338c] = 8'h8d;
s_mem_contents[14'h338d] = 8'h12;
s_mem_contents[14'h338e] = 8'h02;
s_mem_contents[14'h338f] = 8'ha5;
s_mem_contents[14'h3390] = 8'h03;
s_mem_contents[14'h3391] = 8'h20;
s_mem_contents[14'h3392] = 8'h11;
s_mem_contents[14'h3393] = 8'h02;
s_mem_contents[14'h3394] = 8'h08;
s_mem_contents[14'h3395] = 8'hc5;
s_mem_contents[14'h3396] = 8'h05;
s_mem_contents[14'h3397] = 8'hd0;
s_mem_contents[14'h3398] = 8'hfe;
s_mem_contents[14'h3399] = 8'h68;
s_mem_contents[14'h339a] = 8'h29;
s_mem_contents[14'h339b] = 8'hc3;
s_mem_contents[14'h339c] = 8'hc5;
s_mem_contents[14'h339d] = 8'h07;
s_mem_contents[14'h339e] = 8'hd0;
s_mem_contents[14'h339f] = 8'hfe;
s_mem_contents[14'h33a0] = 8'h28;
s_mem_contents[14'h33a1] = 8'h08;
s_mem_contents[14'h33a2] = 8'ha5;
s_mem_contents[14'h33a3] = 8'h08;
s_mem_contents[14'h33a4] = 8'h8d;
s_mem_contents[14'h33a5] = 8'h15;
s_mem_contents[14'h33a6] = 8'h02;
s_mem_contents[14'h33a7] = 8'ha5;
s_mem_contents[14'h33a8] = 8'h03;
s_mem_contents[14'h33a9] = 8'h20;
s_mem_contents[14'h33aa] = 8'h14;
s_mem_contents[14'h33ab] = 8'h02;
s_mem_contents[14'h33ac] = 8'h08;
s_mem_contents[14'h33ad] = 8'hc5;
s_mem_contents[14'h33ae] = 8'h05;
s_mem_contents[14'h33af] = 8'hd0;
s_mem_contents[14'h33b0] = 8'hfe;
s_mem_contents[14'h33b1] = 8'h68;
s_mem_contents[14'h33b2] = 8'h29;
s_mem_contents[14'h33b3] = 8'hc3;
s_mem_contents[14'h33b4] = 8'hc5;
s_mem_contents[14'h33b5] = 8'h07;
s_mem_contents[14'h33b6] = 8'hd0;
s_mem_contents[14'h33b7] = 8'hfe;
s_mem_contents[14'h33b8] = 8'h28;
s_mem_contents[14'h33b9] = 8'h08;
s_mem_contents[14'h33ba] = 8'ha5;
s_mem_contents[14'h33bb] = 8'h03;
s_mem_contents[14'h33bc] = 8'h75;
s_mem_contents[14'h33bd] = 8'h00;
s_mem_contents[14'h33be] = 8'h08;
s_mem_contents[14'h33bf] = 8'hc5;
s_mem_contents[14'h33c0] = 8'h05;
s_mem_contents[14'h33c1] = 8'hd0;
s_mem_contents[14'h33c2] = 8'hfe;
s_mem_contents[14'h33c3] = 8'h68;
s_mem_contents[14'h33c4] = 8'h29;
s_mem_contents[14'h33c5] = 8'hc3;
s_mem_contents[14'h33c6] = 8'hc5;
s_mem_contents[14'h33c7] = 8'h07;
s_mem_contents[14'h33c8] = 8'hd0;
s_mem_contents[14'h33c9] = 8'hfe;
s_mem_contents[14'h33ca] = 8'h28;
s_mem_contents[14'h33cb] = 8'h08;
s_mem_contents[14'h33cc] = 8'ha5;
s_mem_contents[14'h33cd] = 8'h03;
s_mem_contents[14'h33ce] = 8'hf5;
s_mem_contents[14'h33cf] = 8'h04;
s_mem_contents[14'h33d0] = 8'h08;
s_mem_contents[14'h33d1] = 8'hc5;
s_mem_contents[14'h33d2] = 8'h05;
s_mem_contents[14'h33d3] = 8'hd0;
s_mem_contents[14'h33d4] = 8'hfe;
s_mem_contents[14'h33d5] = 8'h68;
s_mem_contents[14'h33d6] = 8'h29;
s_mem_contents[14'h33d7] = 8'hc3;
s_mem_contents[14'h33d8] = 8'hc5;
s_mem_contents[14'h33d9] = 8'h07;
s_mem_contents[14'h33da] = 8'hd0;
s_mem_contents[14'h33db] = 8'hfe;
s_mem_contents[14'h33dc] = 8'h28;
s_mem_contents[14'h33dd] = 8'h08;
s_mem_contents[14'h33de] = 8'ha5;
s_mem_contents[14'h33df] = 8'h03;
s_mem_contents[14'h33e0] = 8'h7d;
s_mem_contents[14'h33e1] = 8'hff;
s_mem_contents[14'h33e2] = 8'h01;
s_mem_contents[14'h33e3] = 8'h08;
s_mem_contents[14'h33e4] = 8'hc5;
s_mem_contents[14'h33e5] = 8'h05;
s_mem_contents[14'h33e6] = 8'hd0;
s_mem_contents[14'h33e7] = 8'hfe;
s_mem_contents[14'h33e8] = 8'h68;
s_mem_contents[14'h33e9] = 8'h29;
s_mem_contents[14'h33ea] = 8'hc3;
s_mem_contents[14'h33eb] = 8'hc5;
s_mem_contents[14'h33ec] = 8'h07;
s_mem_contents[14'h33ed] = 8'hd0;
s_mem_contents[14'h33ee] = 8'hfe;
s_mem_contents[14'h33ef] = 8'h28;
s_mem_contents[14'h33f0] = 8'h08;
s_mem_contents[14'h33f1] = 8'ha5;
s_mem_contents[14'h33f2] = 8'h03;
s_mem_contents[14'h33f3] = 8'hfd;
s_mem_contents[14'h33f4] = 8'h00;
s_mem_contents[14'h33f5] = 8'h02;
s_mem_contents[14'h33f6] = 8'h08;
s_mem_contents[14'h33f7] = 8'hc5;
s_mem_contents[14'h33f8] = 8'h05;
s_mem_contents[14'h33f9] = 8'hd0;
s_mem_contents[14'h33fa] = 8'hfe;
s_mem_contents[14'h33fb] = 8'h68;
s_mem_contents[14'h33fc] = 8'h29;
s_mem_contents[14'h33fd] = 8'hc3;
s_mem_contents[14'h33fe] = 8'hc5;
s_mem_contents[14'h33ff] = 8'h07;
s_mem_contents[14'h3400] = 8'hd0;
s_mem_contents[14'h3401] = 8'hfe;
s_mem_contents[14'h3402] = 8'h28;
s_mem_contents[14'h3403] = 8'h08;
s_mem_contents[14'h3404] = 8'ha5;
s_mem_contents[14'h3405] = 8'h03;
s_mem_contents[14'h3406] = 8'h79;
s_mem_contents[14'h3407] = 8'h04;
s_mem_contents[14'h3408] = 8'h01;
s_mem_contents[14'h3409] = 8'h08;
s_mem_contents[14'h340a] = 8'hc5;
s_mem_contents[14'h340b] = 8'h05;
s_mem_contents[14'h340c] = 8'hd0;
s_mem_contents[14'h340d] = 8'hfe;
s_mem_contents[14'h340e] = 8'h68;
s_mem_contents[14'h340f] = 8'h29;
s_mem_contents[14'h3410] = 8'hc3;
s_mem_contents[14'h3411] = 8'hc5;
s_mem_contents[14'h3412] = 8'h07;
s_mem_contents[14'h3413] = 8'hd0;
s_mem_contents[14'h3414] = 8'hfe;
s_mem_contents[14'h3415] = 8'h28;
s_mem_contents[14'h3416] = 8'h08;
s_mem_contents[14'h3417] = 8'ha5;
s_mem_contents[14'h3418] = 8'h03;
s_mem_contents[14'h3419] = 8'hf9;
s_mem_contents[14'h341a] = 8'h05;
s_mem_contents[14'h341b] = 8'h01;
s_mem_contents[14'h341c] = 8'h08;
s_mem_contents[14'h341d] = 8'hc5;
s_mem_contents[14'h341e] = 8'h05;
s_mem_contents[14'h341f] = 8'hd0;
s_mem_contents[14'h3420] = 8'hfe;
s_mem_contents[14'h3421] = 8'h68;
s_mem_contents[14'h3422] = 8'h29;
s_mem_contents[14'h3423] = 8'hc3;
s_mem_contents[14'h3424] = 8'hc5;
s_mem_contents[14'h3425] = 8'h07;
s_mem_contents[14'h3426] = 8'hd0;
s_mem_contents[14'h3427] = 8'hfe;
s_mem_contents[14'h3428] = 8'h28;
s_mem_contents[14'h3429] = 8'h08;
s_mem_contents[14'h342a] = 8'ha5;
s_mem_contents[14'h342b] = 8'h03;
s_mem_contents[14'h342c] = 8'h61;
s_mem_contents[14'h342d] = 8'h44;
s_mem_contents[14'h342e] = 8'h08;
s_mem_contents[14'h342f] = 8'hc5;
s_mem_contents[14'h3430] = 8'h05;
s_mem_contents[14'h3431] = 8'hd0;
s_mem_contents[14'h3432] = 8'hfe;
s_mem_contents[14'h3433] = 8'h68;
s_mem_contents[14'h3434] = 8'h29;
s_mem_contents[14'h3435] = 8'hc3;
s_mem_contents[14'h3436] = 8'hc5;
s_mem_contents[14'h3437] = 8'h07;
s_mem_contents[14'h3438] = 8'hd0;
s_mem_contents[14'h3439] = 8'hfe;
s_mem_contents[14'h343a] = 8'h28;
s_mem_contents[14'h343b] = 8'h08;
s_mem_contents[14'h343c] = 8'ha5;
s_mem_contents[14'h343d] = 8'h03;
s_mem_contents[14'h343e] = 8'he1;
s_mem_contents[14'h343f] = 8'h46;
s_mem_contents[14'h3440] = 8'h08;
s_mem_contents[14'h3441] = 8'hc5;
s_mem_contents[14'h3442] = 8'h05;
s_mem_contents[14'h3443] = 8'hd0;
s_mem_contents[14'h3444] = 8'hfe;
s_mem_contents[14'h3445] = 8'h68;
s_mem_contents[14'h3446] = 8'h29;
s_mem_contents[14'h3447] = 8'hc3;
s_mem_contents[14'h3448] = 8'hc5;
s_mem_contents[14'h3449] = 8'h07;
s_mem_contents[14'h344a] = 8'hd0;
s_mem_contents[14'h344b] = 8'hfe;
s_mem_contents[14'h344c] = 8'h28;
s_mem_contents[14'h344d] = 8'h08;
s_mem_contents[14'h344e] = 8'ha5;
s_mem_contents[14'h344f] = 8'h03;
s_mem_contents[14'h3450] = 8'h71;
s_mem_contents[14'h3451] = 8'h4c;
s_mem_contents[14'h3452] = 8'h08;
s_mem_contents[14'h3453] = 8'hc5;
s_mem_contents[14'h3454] = 8'h05;
s_mem_contents[14'h3455] = 8'hd0;
s_mem_contents[14'h3456] = 8'hfe;
s_mem_contents[14'h3457] = 8'h68;
s_mem_contents[14'h3458] = 8'h29;
s_mem_contents[14'h3459] = 8'hc3;
s_mem_contents[14'h345a] = 8'hc5;
s_mem_contents[14'h345b] = 8'h07;
s_mem_contents[14'h345c] = 8'hd0;
s_mem_contents[14'h345d] = 8'hfe;
s_mem_contents[14'h345e] = 8'h28;
s_mem_contents[14'h345f] = 8'h08;
s_mem_contents[14'h3460] = 8'ha5;
s_mem_contents[14'h3461] = 8'h03;
s_mem_contents[14'h3462] = 8'hf1;
s_mem_contents[14'h3463] = 8'h4e;
s_mem_contents[14'h3464] = 8'h08;
s_mem_contents[14'h3465] = 8'hc5;
s_mem_contents[14'h3466] = 8'h05;
s_mem_contents[14'h3467] = 8'hd0;
s_mem_contents[14'h3468] = 8'hfe;
s_mem_contents[14'h3469] = 8'h68;
s_mem_contents[14'h346a] = 8'h29;
s_mem_contents[14'h346b] = 8'hc3;
s_mem_contents[14'h346c] = 8'hc5;
s_mem_contents[14'h346d] = 8'h07;
s_mem_contents[14'h346e] = 8'hd0;
s_mem_contents[14'h346f] = 8'hfe;
s_mem_contents[14'h3470] = 8'h28;
s_mem_contents[14'h3471] = 8'h60;
s_mem_contents[14'h3472] = 8'h88;
s_mem_contents[14'h3473] = 8'h88;
s_mem_contents[14'h3474] = 8'h08;
s_mem_contents[14'h3475] = 8'h88;
s_mem_contents[14'h3476] = 8'h88;
s_mem_contents[14'h3477] = 8'h88;
s_mem_contents[14'h3478] = 8'h28;
s_mem_contents[14'h3479] = 8'hb0;
s_mem_contents[14'h347a] = 8'hfe;
s_mem_contents[14'h347b] = 8'h70;
s_mem_contents[14'h347c] = 8'hfe;
s_mem_contents[14'h347d] = 8'h30;
s_mem_contents[14'h347e] = 8'hfe;
s_mem_contents[14'h347f] = 8'hf0;
s_mem_contents[14'h3480] = 8'hfe;
s_mem_contents[14'h3481] = 8'hc9;
s_mem_contents[14'h3482] = 8'h46;
s_mem_contents[14'h3483] = 8'hd0;
s_mem_contents[14'h3484] = 8'hfe;
s_mem_contents[14'h3485] = 8'he0;
s_mem_contents[14'h3486] = 8'h41;
s_mem_contents[14'h3487] = 8'hd0;
s_mem_contents[14'h3488] = 8'hfe;
s_mem_contents[14'h3489] = 8'hc0;
s_mem_contents[14'h348a] = 8'h4f;
s_mem_contents[14'h348b] = 8'hd0;
s_mem_contents[14'h348c] = 8'hfe;
s_mem_contents[14'h348d] = 8'h48;
s_mem_contents[14'h348e] = 8'h8a;
s_mem_contents[14'h348f] = 8'h48;
s_mem_contents[14'h3490] = 8'hba;
s_mem_contents[14'h3491] = 8'he0;
s_mem_contents[14'h3492] = 8'hfd;
s_mem_contents[14'h3493] = 8'hd0;
s_mem_contents[14'h3494] = 8'hfe;
s_mem_contents[14'h3495] = 8'h68;
s_mem_contents[14'h3496] = 8'haa;
s_mem_contents[14'h3497] = 8'ha9;
s_mem_contents[14'h3498] = 8'hff;
s_mem_contents[14'h3499] = 8'h48;
s_mem_contents[14'h349a] = 8'h28;
s_mem_contents[14'h349b] = 8'h68;
s_mem_contents[14'h349c] = 8'he8;
s_mem_contents[14'h349d] = 8'h49;
s_mem_contents[14'h349e] = 8'haa;
s_mem_contents[14'h349f] = 8'h4c;
s_mem_contents[14'h34a0] = 8'h0f;
s_mem_contents[14'h34a1] = 8'h09;
s_mem_contents[14'h34a2] = 8'hab;
s_mem_contents[14'h34a3] = 8'h34;
s_mem_contents[14'h34a4] = 8'h64;
s_mem_contents[14'h34a5] = 8'h09;
s_mem_contents[14'h34a6] = 8'h4c;
s_mem_contents[14'h34a7] = 8'ha6;
s_mem_contents[14'h34a8] = 8'h34;
s_mem_contents[14'h34a9] = 8'h88;
s_mem_contents[14'h34aa] = 8'h88;
s_mem_contents[14'h34ab] = 8'h08;
s_mem_contents[14'h34ac] = 8'h88;
s_mem_contents[14'h34ad] = 8'h88;
s_mem_contents[14'h34ae] = 8'h88;
s_mem_contents[14'h34af] = 8'h28;
s_mem_contents[14'h34b0] = 8'hb0;
s_mem_contents[14'h34b1] = 8'hfe;
s_mem_contents[14'h34b2] = 8'h70;
s_mem_contents[14'h34b3] = 8'hfe;
s_mem_contents[14'h34b4] = 8'h30;
s_mem_contents[14'h34b5] = 8'hfe;
s_mem_contents[14'h34b6] = 8'hf0;
s_mem_contents[14'h34b7] = 8'hfe;
s_mem_contents[14'h34b8] = 8'hc9;
s_mem_contents[14'h34b9] = 8'h49;
s_mem_contents[14'h34ba] = 8'hd0;
s_mem_contents[14'h34bb] = 8'hfe;
s_mem_contents[14'h34bc] = 8'he0;
s_mem_contents[14'h34bd] = 8'h4e;
s_mem_contents[14'h34be] = 8'hd0;
s_mem_contents[14'h34bf] = 8'hfe;
s_mem_contents[14'h34c0] = 8'hc0;
s_mem_contents[14'h34c1] = 8'h41;
s_mem_contents[14'h34c2] = 8'hd0;
s_mem_contents[14'h34c3] = 8'hfe;
s_mem_contents[14'h34c4] = 8'h48;
s_mem_contents[14'h34c5] = 8'h8a;
s_mem_contents[14'h34c6] = 8'h48;
s_mem_contents[14'h34c7] = 8'hba;
s_mem_contents[14'h34c8] = 8'he0;
s_mem_contents[14'h34c9] = 8'hfd;
s_mem_contents[14'h34ca] = 8'hd0;
s_mem_contents[14'h34cb] = 8'hfe;
s_mem_contents[14'h34cc] = 8'h68;
s_mem_contents[14'h34cd] = 8'haa;
s_mem_contents[14'h34ce] = 8'ha9;
s_mem_contents[14'h34cf] = 8'hff;
s_mem_contents[14'h34d0] = 8'h48;
s_mem_contents[14'h34d1] = 8'h28;
s_mem_contents[14'h34d2] = 8'h68;
s_mem_contents[14'h34d3] = 8'he8;
s_mem_contents[14'h34d4] = 8'h49;
s_mem_contents[14'h34d5] = 8'haa;
s_mem_contents[14'h34d6] = 8'h6c;
s_mem_contents[14'h34d7] = 8'ha4;
s_mem_contents[14'h34d8] = 8'h34;
s_mem_contents[14'h34d9] = 8'h4c;
s_mem_contents[14'h34da] = 8'hd9;
s_mem_contents[14'h34db] = 8'h34;
s_mem_contents[14'h34dc] = 8'h4c;
s_mem_contents[14'h34dd] = 8'h00;
s_mem_contents[14'h34de] = 8'h04;
s_mem_contents[14'h34df] = 8'h88;
s_mem_contents[14'h34e0] = 8'h88;
s_mem_contents[14'h34e1] = 8'h08;
s_mem_contents[14'h34e2] = 8'h88;
s_mem_contents[14'h34e3] = 8'h88;
s_mem_contents[14'h34e4] = 8'h88;
s_mem_contents[14'h34e5] = 8'h28;
s_mem_contents[14'h34e6] = 8'hb0;
s_mem_contents[14'h34e7] = 8'hfe;
s_mem_contents[14'h34e8] = 8'h70;
s_mem_contents[14'h34e9] = 8'hfe;
s_mem_contents[14'h34ea] = 8'h30;
s_mem_contents[14'h34eb] = 8'hfe;
s_mem_contents[14'h34ec] = 8'hf0;
s_mem_contents[14'h34ed] = 8'hfe;
s_mem_contents[14'h34ee] = 8'hc9;
s_mem_contents[14'h34ef] = 8'h4a;
s_mem_contents[14'h34f0] = 8'hd0;
s_mem_contents[14'h34f1] = 8'hfe;
s_mem_contents[14'h34f2] = 8'he0;
s_mem_contents[14'h34f3] = 8'h53;
s_mem_contents[14'h34f4] = 8'hd0;
s_mem_contents[14'h34f5] = 8'hfe;
s_mem_contents[14'h34f6] = 8'hc0;
s_mem_contents[14'h34f7] = 8'h4f;
s_mem_contents[14'h34f8] = 8'hd0;
s_mem_contents[14'h34f9] = 8'hfe;
s_mem_contents[14'h34fa] = 8'h48;
s_mem_contents[14'h34fb] = 8'h8a;
s_mem_contents[14'h34fc] = 8'h48;
s_mem_contents[14'h34fd] = 8'hba;
s_mem_contents[14'h34fe] = 8'he0;
s_mem_contents[14'h34ff] = 8'hfb;
s_mem_contents[14'h3500] = 8'hd0;
s_mem_contents[14'h3501] = 8'hfe;
s_mem_contents[14'h3502] = 8'had;
s_mem_contents[14'h3503] = 8'hff;
s_mem_contents[14'h3504] = 8'h01;
s_mem_contents[14'h3505] = 8'hc9;
s_mem_contents[14'h3506] = 8'h09;
s_mem_contents[14'h3507] = 8'hd0;
s_mem_contents[14'h3508] = 8'hfe;
s_mem_contents[14'h3509] = 8'had;
s_mem_contents[14'h350a] = 8'hfe;
s_mem_contents[14'h350b] = 8'h01;
s_mem_contents[14'h350c] = 8'hc9;
s_mem_contents[14'h350d] = 8'h9a;
s_mem_contents[14'h350e] = 8'hd0;
s_mem_contents[14'h350f] = 8'hfe;
s_mem_contents[14'h3510] = 8'ha9;
s_mem_contents[14'h3511] = 8'hff;
s_mem_contents[14'h3512] = 8'h48;
s_mem_contents[14'h3513] = 8'h28;
s_mem_contents[14'h3514] = 8'h68;
s_mem_contents[14'h3515] = 8'haa;
s_mem_contents[14'h3516] = 8'h68;
s_mem_contents[14'h3517] = 8'he8;
s_mem_contents[14'h3518] = 8'h49;
s_mem_contents[14'h3519] = 8'haa;
s_mem_contents[14'h351a] = 8'h60;
s_mem_contents[14'h351b] = 8'h4c;
s_mem_contents[14'h351c] = 8'h1b;
s_mem_contents[14'h351d] = 8'h35;
s_mem_contents[14'h351e] = 8'h4c;
s_mem_contents[14'h351f] = 8'h00;
s_mem_contents[14'h3520] = 8'h04;
s_mem_contents[14'h3521] = 8'h4c;
s_mem_contents[14'h3522] = 8'h21;
s_mem_contents[14'h3523] = 8'h35;
s_mem_contents[14'h3524] = 8'h4c;
s_mem_contents[14'h3525] = 8'h00;
s_mem_contents[14'h3526] = 8'h04;
s_mem_contents[14'h3527] = 8'h4c;
s_mem_contents[14'h3528] = 8'h27;
s_mem_contents[14'h3529] = 8'h35;
s_mem_contents[14'h352a] = 8'h4c;
s_mem_contents[14'h352b] = 8'h00;
s_mem_contents[14'h352c] = 8'h04;
s_mem_contents[14'h352d] = 8'h88;
s_mem_contents[14'h352e] = 8'h88;

`endif

  end

  always @(posedge CLK) begin
    if (WE)
      s_mem_contents[Address[13:0]] <= DataIn;
    else
      DataOut <= s_mem_contents[Address[13:0]];
  end

endmodule
