/*module fsm(
  input AB,
  input ACI,
  input CLK,
  input[1:0] GR,
  input ID,
  input[2:0] OPC,
  input R,
  input XY,
  output ACO,
  output ADR,
  output ALU,
  output[5:0] AOP,
  output INC,
  output LCO,
  output MHI,
  output MLO,
  output PRV,
  output rX,
  output rY,
  output wA,
  output wL,
  output wO,
  output wX,
  output wY
);

endmodule
*/
