module bitmap(
  input CLK,
  input WE,
  input[13:0] Address,
  input[7:0] DataIn,
  output reg[7:0] DataOut
);

  // 320x200 / 8 = 8000
  // 16000 gives 2 monochrome images
  reg [7:0] memory[15999:0];
  parameter base = 8000;

  integer i,j;
  initial begin
/*
    for (i=0;i<40;i=i+1) begin
      for (j=0;j<200;j=j+1) begin
        if (j % 8 && (i == 0 || i == 39))
          memory[base+j*40+i] = 8'b01111111;
        if (j > 4-4 && j < 4+4)
          memory[base+j*40+i] = 8'b01111111;
        if (j > 92-4 && j < 92+4) begin
          memory[base+j*40+i] = 8'b01111111;
        end
        if (j > 100-4 && j < 100+4) begin
          memory[base+j*40+i] = 8'b01111111;
        end
        if (j > 108-4 && j < 108+4) begin
          memory[base+j*40+i] = 8'b01111111;
        end
        if (j > 196-4 && j < 196+4)
          memory[base+j*40+i] = 8'b01111111;
      end
    end
*/
///*
memory[0]=8'b11111111;
memory[1]=8'b11111111;
memory[2]=8'b11111111;
memory[3]=8'b11111111;
memory[4]=8'b11111111;
memory[5]=8'b11111111;
memory[6]=8'b11111111;
memory[7]=8'b11111111;
memory[8]=8'b11111111;
memory[9]=8'b11111111;
memory[10]=8'b11111111;
memory[11]=8'b11111111;
memory[12]=8'b11111111;
memory[13]=8'b11111111;
memory[14]=8'b11111111;
memory[15]=8'b11111111;
memory[16]=8'b11111111;
memory[17]=8'b11111111;
memory[18]=8'b11111111;
memory[19]=8'b11111111;
memory[20]=8'b11111111;
memory[21]=8'b11111111;
memory[22]=8'b11111111;
memory[23]=8'b11111111;
memory[24]=8'b11111111;
memory[25]=8'b11111111;
memory[26]=8'b11111111;
memory[27]=8'b11111111;
memory[28]=8'b11111111;
memory[29]=8'b11111111;
memory[30]=8'b11111111;
memory[31]=8'b11111111;
memory[32]=8'b11111111;
memory[33]=8'b11111111;
memory[34]=8'b11111111;
memory[35]=8'b11111111;
memory[36]=8'b11111111;
memory[37]=8'b11111111;
memory[38]=8'b11111111;
memory[39]=8'b11111111;
memory[40]=8'b11111111;
memory[41]=8'b11111111;
memory[42]=8'b11111111;
memory[43]=8'b11111111;
memory[44]=8'b11111111;
memory[45]=8'b11111111;
memory[46]=8'b11111111;
memory[47]=8'b11111111;
memory[48]=8'b11111111;
memory[49]=8'b11111111;
memory[50]=8'b11111111;
memory[51]=8'b11111111;
memory[52]=8'b11111111;
memory[53]=8'b11111111;
memory[54]=8'b11111111;
memory[55]=8'b11111111;
memory[56]=8'b11111111;
memory[57]=8'b11111111;
memory[58]=8'b11111111;
memory[59]=8'b11111111;
memory[60]=8'b11111111;
memory[61]=8'b11111111;
memory[62]=8'b11111111;
memory[63]=8'b11111111;
memory[64]=8'b11111111;
memory[65]=8'b11111111;
memory[66]=8'b11111111;
memory[67]=8'b11111111;
memory[68]=8'b11111111;
memory[69]=8'b11111111;
memory[70]=8'b11111111;
memory[71]=8'b11111111;
memory[72]=8'b11111111;
memory[73]=8'b11111111;
memory[74]=8'b11111111;
memory[75]=8'b11111111;
memory[76]=8'b11111111;
memory[77]=8'b11111111;
memory[78]=8'b11111111;
memory[79]=8'b11111111;
memory[80]=8'b11111111;
memory[81]=8'b11111111;
memory[82]=8'b11111111;
memory[83]=8'b11111111;
memory[84]=8'b11111111;
memory[85]=8'b11111111;
memory[86]=8'b11111111;
memory[87]=8'b11111111;
memory[88]=8'b11111111;
memory[89]=8'b11111111;
memory[90]=8'b11111111;
memory[91]=8'b11111111;
memory[92]=8'b11111111;
memory[93]=8'b11111111;
memory[94]=8'b11111111;
memory[95]=8'b11111111;
memory[96]=8'b11111111;
memory[97]=8'b11111111;
memory[98]=8'b11111111;
memory[99]=8'b11111111;
memory[100]=8'b11111111;
memory[101]=8'b11111111;
memory[102]=8'b11111111;
memory[103]=8'b11111111;
memory[104]=8'b11111111;
memory[105]=8'b11111111;
memory[106]=8'b11111111;
memory[107]=8'b11111111;
memory[108]=8'b11111111;
memory[109]=8'b11111111;
memory[110]=8'b11111111;
memory[111]=8'b11111111;
memory[112]=8'b11111111;
memory[113]=8'b11111111;
memory[114]=8'b11111111;
memory[115]=8'b11111111;
memory[116]=8'b11111111;
memory[117]=8'b11111111;
memory[118]=8'b11111111;
memory[119]=8'b11111111;
memory[120]=8'b11111111;
memory[121]=8'b11111111;
memory[122]=8'b11111111;
memory[123]=8'b11111111;
memory[124]=8'b11111111;
memory[125]=8'b11111111;
memory[126]=8'b11111111;
memory[127]=8'b11111111;
memory[128]=8'b11111111;
memory[129]=8'b11111111;
memory[130]=8'b11111111;
memory[131]=8'b11111111;
memory[132]=8'b11111111;
memory[133]=8'b11111111;
memory[134]=8'b11111111;
memory[135]=8'b11111111;
memory[136]=8'b11111111;
memory[137]=8'b11111111;
memory[138]=8'b11111111;
memory[139]=8'b11111111;
memory[140]=8'b11111111;
memory[141]=8'b11111111;
memory[142]=8'b11111111;
memory[143]=8'b11111111;
memory[144]=8'b11111111;
memory[145]=8'b11111111;
memory[146]=8'b11111111;
memory[147]=8'b11111111;
memory[148]=8'b11111111;
memory[149]=8'b11111111;
memory[150]=8'b11111111;
memory[151]=8'b11111111;
memory[152]=8'b11111111;
memory[153]=8'b11111111;
memory[154]=8'b11111111;
memory[155]=8'b11111111;
memory[156]=8'b11111111;
memory[157]=8'b11111111;
memory[158]=8'b11111111;
memory[159]=8'b11111111;
memory[160]=8'b11111111;
memory[161]=8'b11111111;
memory[162]=8'b11111111;
memory[163]=8'b11111111;
memory[164]=8'b11111111;
memory[165]=8'b11111111;
memory[166]=8'b11111111;
memory[167]=8'b11111111;
memory[168]=8'b11111111;
memory[169]=8'b11111111;
memory[170]=8'b11111111;
memory[171]=8'b11111111;
memory[172]=8'b11111111;
memory[173]=8'b11111111;
memory[174]=8'b11111111;
memory[175]=8'b11111111;
memory[176]=8'b11111111;
memory[177]=8'b11111111;
memory[178]=8'b11111111;
memory[179]=8'b11111111;
memory[180]=8'b11111111;
memory[181]=8'b11111111;
memory[182]=8'b11111111;
memory[183]=8'b11111111;
memory[184]=8'b11111111;
memory[185]=8'b11111111;
memory[186]=8'b11111111;
memory[187]=8'b11111111;
memory[188]=8'b11111111;
memory[189]=8'b11111111;
memory[190]=8'b11111111;
memory[191]=8'b11111111;
memory[192]=8'b11111111;
memory[193]=8'b11111111;
memory[194]=8'b11111111;
memory[195]=8'b11111111;
memory[196]=8'b11111111;
memory[197]=8'b11111111;
memory[198]=8'b11111111;
memory[199]=8'b11111111;
memory[200]=8'b11111111;
memory[201]=8'b11111111;
memory[202]=8'b11111111;
memory[203]=8'b11111111;
memory[204]=8'b11111111;
memory[205]=8'b11111111;
memory[206]=8'b11111111;
memory[207]=8'b11111111;
memory[208]=8'b11111111;
memory[209]=8'b11111111;
memory[210]=8'b11111111;
memory[211]=8'b11111111;
memory[212]=8'b11111111;
memory[213]=8'b11111111;
memory[214]=8'b11111111;
memory[215]=8'b11111111;
memory[216]=8'b11111111;
memory[217]=8'b11111111;
memory[218]=8'b11111111;
memory[219]=8'b11111111;
memory[220]=8'b11111111;
memory[221]=8'b11111111;
memory[222]=8'b11111111;
memory[223]=8'b11111111;
memory[224]=8'b11111111;
memory[225]=8'b11111111;
memory[226]=8'b11111111;
memory[227]=8'b11111111;
memory[228]=8'b11111111;
memory[229]=8'b11111111;
memory[230]=8'b11111111;
memory[231]=8'b11111111;
memory[232]=8'b11111111;
memory[233]=8'b11111111;
memory[234]=8'b11111111;
memory[235]=8'b11111111;
memory[236]=8'b11111111;
memory[237]=8'b11111111;
memory[238]=8'b11111111;
memory[239]=8'b11111111;
memory[240]=8'b11111111;
memory[241]=8'b11111111;
memory[242]=8'b11111111;
memory[243]=8'b11111111;
memory[244]=8'b11111111;
memory[245]=8'b11111111;
memory[246]=8'b11111111;
memory[247]=8'b11111111;
memory[248]=8'b11111111;
memory[249]=8'b11111111;
memory[250]=8'b11111111;
memory[251]=8'b11111111;
memory[252]=8'b11111111;
memory[253]=8'b11111111;
memory[254]=8'b11111111;
memory[255]=8'b11111111;
memory[256]=8'b11111111;
memory[257]=8'b11111111;
memory[258]=8'b11111111;
memory[259]=8'b11111111;
memory[260]=8'b11111111;
memory[261]=8'b11111111;
memory[262]=8'b11111111;
memory[263]=8'b11111111;
memory[264]=8'b11111111;
memory[265]=8'b11111111;
memory[266]=8'b11111111;
memory[267]=8'b11111111;
memory[268]=8'b11111111;
memory[269]=8'b11111111;
memory[270]=8'b11111111;
memory[271]=8'b11111111;
memory[272]=8'b11111111;
memory[273]=8'b11111111;
memory[274]=8'b11111111;
memory[275]=8'b11111111;
memory[276]=8'b11111111;
memory[277]=8'b11111111;
memory[278]=8'b11111111;
memory[279]=8'b11111111;
memory[280]=8'b11111111;
memory[281]=8'b11111111;
memory[282]=8'b11111111;
memory[283]=8'b11111111;
memory[284]=8'b11111111;
memory[285]=8'b11111111;
memory[286]=8'b11111111;
memory[287]=8'b11111111;
memory[288]=8'b11111111;
memory[289]=8'b11111111;
memory[290]=8'b11111111;
memory[291]=8'b11111111;
memory[292]=8'b11111111;
memory[293]=8'b11111111;
memory[294]=8'b11111111;
memory[295]=8'b11111111;
memory[296]=8'b11111111;
memory[297]=8'b11111111;
memory[298]=8'b11111111;
memory[299]=8'b11111111;
memory[300]=8'b11111111;
memory[301]=8'b11111111;
memory[302]=8'b11111111;
memory[303]=8'b11111111;
memory[304]=8'b11111111;
memory[305]=8'b11111111;
memory[306]=8'b11111111;
memory[307]=8'b11111111;
memory[308]=8'b11111111;
memory[309]=8'b11111111;
memory[310]=8'b11111111;
memory[311]=8'b11111111;
memory[312]=8'b11111111;
memory[313]=8'b11111111;
memory[314]=8'b11111111;
memory[315]=8'b11111111;
memory[316]=8'b11111111;
memory[317]=8'b11111111;
memory[318]=8'b11111111;
memory[319]=8'b11111111;
memory[320]=8'b11111111;
memory[321]=8'b11111111;
memory[322]=8'b11111111;
memory[323]=8'b11111111;
memory[324]=8'b11111111;
memory[325]=8'b11111111;
memory[326]=8'b11111111;
memory[327]=8'b11111111;
memory[328]=8'b11111111;
memory[329]=8'b11111111;
memory[330]=8'b11111111;
memory[331]=8'b11111111;
memory[332]=8'b11111111;
memory[333]=8'b11111111;
memory[334]=8'b11111111;
memory[335]=8'b11111111;
memory[336]=8'b11111111;
memory[337]=8'b11111111;
memory[338]=8'b11111111;
memory[339]=8'b11111111;
memory[340]=8'b11111111;
memory[341]=8'b11111111;
memory[342]=8'b11111111;
memory[343]=8'b11111111;
memory[344]=8'b11111111;
memory[345]=8'b11111111;
memory[346]=8'b11111111;
memory[347]=8'b11111111;
memory[348]=8'b11111111;
memory[349]=8'b11111111;
memory[350]=8'b11111111;
memory[351]=8'b11111111;
memory[352]=8'b11111111;
memory[353]=8'b11111111;
memory[354]=8'b11111111;
memory[355]=8'b11111111;
memory[356]=8'b11111111;
memory[357]=8'b11111111;
memory[358]=8'b11111111;
memory[359]=8'b11111111;
memory[360]=8'b11111111;
memory[361]=8'b11111111;
memory[362]=8'b11111111;
memory[363]=8'b11111111;
memory[364]=8'b11111111;
memory[365]=8'b11111111;
memory[366]=8'b11111111;
memory[367]=8'b11111111;
memory[368]=8'b11111111;
memory[369]=8'b11111111;
memory[370]=8'b11111111;
memory[371]=8'b11111111;
memory[372]=8'b11111111;
memory[373]=8'b11111111;
memory[374]=8'b11111111;
memory[375]=8'b11111111;
memory[376]=8'b11111111;
memory[377]=8'b11111111;
memory[378]=8'b11111111;
memory[379]=8'b11111111;
memory[380]=8'b11111111;
memory[381]=8'b11111111;
memory[382]=8'b11111111;
memory[383]=8'b11111111;
memory[384]=8'b11111111;
memory[385]=8'b11111111;
memory[386]=8'b11111111;
memory[387]=8'b11111111;
memory[388]=8'b11111111;
memory[389]=8'b11111111;
memory[390]=8'b11111111;
memory[391]=8'b11111111;
memory[392]=8'b11111111;
memory[393]=8'b11111111;
memory[394]=8'b11111111;
memory[395]=8'b11111111;
memory[396]=8'b11111111;
memory[397]=8'b11111111;
memory[398]=8'b11111111;
memory[399]=8'b11111111;
memory[400]=8'b11111111;
memory[401]=8'b11111111;
memory[402]=8'b11111111;
memory[403]=8'b11111111;
memory[404]=8'b11111111;
memory[405]=8'b11111111;
memory[406]=8'b11111111;
memory[407]=8'b11111111;
memory[408]=8'b11111111;
memory[409]=8'b11111111;
memory[410]=8'b11111111;
memory[411]=8'b11111111;
memory[412]=8'b11111111;
memory[413]=8'b11111111;
memory[414]=8'b11111111;
memory[415]=8'b11111111;
memory[416]=8'b11111111;
memory[417]=8'b11111111;
memory[418]=8'b11111111;
memory[419]=8'b11111111;
memory[420]=8'b11111111;
memory[421]=8'b11111000;
memory[422]=8'b00001111;
memory[423]=8'b11111111;
memory[424]=8'b11111111;
memory[425]=8'b11111111;
memory[426]=8'b11111111;
memory[427]=8'b11111111;
memory[428]=8'b11111111;
memory[429]=8'b11111111;
memory[430]=8'b11111111;
memory[431]=8'b11111111;
memory[432]=8'b11111111;
memory[433]=8'b11111111;
memory[434]=8'b11111111;
memory[435]=8'b11111111;
memory[436]=8'b11111111;
memory[437]=8'b11111111;
memory[438]=8'b11111111;
memory[439]=8'b11111111;
memory[440]=8'b11111111;
memory[441]=8'b11111111;
memory[442]=8'b11111111;
memory[443]=8'b11111111;
memory[444]=8'b11111111;
memory[445]=8'b11111111;
memory[446]=8'b11111111;
memory[447]=8'b11111111;
memory[448]=8'b11111111;
memory[449]=8'b11111111;
memory[450]=8'b11111111;
memory[451]=8'b11111111;
memory[452]=8'b11111111;
memory[453]=8'b11111111;
memory[454]=8'b11111111;
memory[455]=8'b11111111;
memory[456]=8'b11111111;
memory[457]=8'b11111111;
memory[458]=8'b11111111;
memory[459]=8'b11111111;
memory[460]=8'b11111111;
memory[461]=8'b10000000;
memory[462]=8'b00000001;
memory[463]=8'b11111111;
memory[464]=8'b11111111;
memory[465]=8'b11111111;
memory[466]=8'b11111111;
memory[467]=8'b11111111;
memory[468]=8'b11111111;
memory[469]=8'b11111111;
memory[470]=8'b11111111;
memory[471]=8'b11111111;
memory[472]=8'b11111111;
memory[473]=8'b11111111;
memory[474]=8'b11111111;
memory[475]=8'b11111111;
memory[476]=8'b11111111;
memory[477]=8'b11111111;
memory[478]=8'b11111111;
memory[479]=8'b11111111;
memory[480]=8'b11111111;
memory[481]=8'b11111111;
memory[482]=8'b11111111;
memory[483]=8'b11111111;
memory[484]=8'b11111111;
memory[485]=8'b11111111;
memory[486]=8'b11111111;
memory[487]=8'b11111111;
memory[488]=8'b11111111;
memory[489]=8'b11111111;
memory[490]=8'b11111111;
memory[491]=8'b11111111;
memory[492]=8'b11111111;
memory[493]=8'b11111111;
memory[494]=8'b11111111;
memory[495]=8'b11111111;
memory[496]=8'b11111111;
memory[497]=8'b11111111;
memory[498]=8'b11111111;
memory[499]=8'b11111111;
memory[500]=8'b11111110;
memory[501]=8'b00000000;
memory[502]=8'b00000000;
memory[503]=8'b01111111;
memory[504]=8'b11111111;
memory[505]=8'b11111111;
memory[506]=8'b11111111;
memory[507]=8'b11111111;
memory[508]=8'b11111111;
memory[509]=8'b11111111;
memory[510]=8'b11111111;
memory[511]=8'b11111111;
memory[512]=8'b11111111;
memory[513]=8'b11111111;
memory[514]=8'b11111111;
memory[515]=8'b11111111;
memory[516]=8'b11111111;
memory[517]=8'b11111111;
memory[518]=8'b11111111;
memory[519]=8'b11111111;
memory[520]=8'b11111111;
memory[521]=8'b11111111;
memory[522]=8'b11111111;
memory[523]=8'b11111111;
memory[524]=8'b11111111;
memory[525]=8'b11111111;
memory[526]=8'b11111111;
memory[527]=8'b11111111;
memory[528]=8'b11111111;
memory[529]=8'b11111111;
memory[530]=8'b11111111;
memory[531]=8'b11111111;
memory[532]=8'b11111111;
memory[533]=8'b11111111;
memory[534]=8'b11111111;
memory[535]=8'b11111111;
memory[536]=8'b11111111;
memory[537]=8'b11111111;
memory[538]=8'b11111111;
memory[539]=8'b11111111;
memory[540]=8'b11111100;
memory[541]=8'b00000000;
memory[542]=8'b00000000;
memory[543]=8'b00111111;
memory[544]=8'b11111111;
memory[545]=8'b11111111;
memory[546]=8'b11111111;
memory[547]=8'b11111111;
memory[548]=8'b11111111;
memory[549]=8'b11111111;
memory[550]=8'b11111111;
memory[551]=8'b11111111;
memory[552]=8'b11111111;
memory[553]=8'b11111111;
memory[554]=8'b11111111;
memory[555]=8'b11111111;
memory[556]=8'b11111111;
memory[557]=8'b11111111;
memory[558]=8'b11111111;
memory[559]=8'b11111111;
memory[560]=8'b11111111;
memory[561]=8'b11111111;
memory[562]=8'b11111111;
memory[563]=8'b11111111;
memory[564]=8'b11111111;
memory[565]=8'b11111111;
memory[566]=8'b11111111;
memory[567]=8'b11111111;
memory[568]=8'b11111111;
memory[569]=8'b11111111;
memory[570]=8'b11111111;
memory[571]=8'b11111111;
memory[572]=8'b11111111;
memory[573]=8'b11111111;
memory[574]=8'b11111111;
memory[575]=8'b11111111;
memory[576]=8'b11111111;
memory[577]=8'b11111111;
memory[578]=8'b11111111;
memory[579]=8'b11111111;
memory[580]=8'b11111000;
memory[581]=8'b00000000;
memory[582]=8'b00000000;
memory[583]=8'b00001111;
memory[584]=8'b11111111;
memory[585]=8'b11111111;
memory[586]=8'b11111111;
memory[587]=8'b11111111;
memory[588]=8'b11111111;
memory[589]=8'b11111111;
memory[590]=8'b11001111;
memory[591]=8'b11111111;
memory[592]=8'b11111111;
memory[593]=8'b11111111;
memory[594]=8'b11111111;
memory[595]=8'b11111111;
memory[596]=8'b11111111;
memory[597]=8'b11111111;
memory[598]=8'b11111111;
memory[599]=8'b11111111;
memory[600]=8'b11111111;
memory[601]=8'b11111111;
memory[602]=8'b11111111;
memory[603]=8'b11111111;
memory[604]=8'b11111111;
memory[605]=8'b11111111;
memory[606]=8'b11111111;
memory[607]=8'b11111111;
memory[608]=8'b11111111;
memory[609]=8'b11111111;
memory[610]=8'b11111111;
memory[611]=8'b11111111;
memory[612]=8'b11111111;
memory[613]=8'b11111111;
memory[614]=8'b11111111;
memory[615]=8'b11111111;
memory[616]=8'b11111111;
memory[617]=8'b11111111;
memory[618]=8'b11111111;
memory[619]=8'b11111111;
memory[620]=8'b11110000;
memory[621]=8'b00000000;
memory[622]=8'b00000000;
memory[623]=8'b00001111;
memory[624]=8'b11111111;
memory[625]=8'b11111111;
memory[626]=8'b11111111;
memory[627]=8'b11111111;
memory[628]=8'b11111111;
memory[629]=8'b11111111;
memory[630]=8'b10000111;
memory[631]=8'b11111111;
memory[632]=8'b11111111;
memory[633]=8'b11111111;
memory[634]=8'b11111111;
memory[635]=8'b11111111;
memory[636]=8'b11111111;
memory[637]=8'b11111111;
memory[638]=8'b11111111;
memory[639]=8'b11111111;
memory[640]=8'b11111111;
memory[641]=8'b11111111;
memory[642]=8'b11111111;
memory[643]=8'b11111111;
memory[644]=8'b11111111;
memory[645]=8'b11111111;
memory[646]=8'b11111111;
memory[647]=8'b11111111;
memory[648]=8'b11111111;
memory[649]=8'b11111111;
memory[650]=8'b11111111;
memory[651]=8'b11111111;
memory[652]=8'b11111111;
memory[653]=8'b11111111;
memory[654]=8'b11111111;
memory[655]=8'b11111111;
memory[656]=8'b11111111;
memory[657]=8'b11111111;
memory[658]=8'b11111111;
memory[659]=8'b11111111;
memory[660]=8'b11110000;
memory[661]=8'b00000000;
memory[662]=8'b00000000;
memory[663]=8'b00000111;
memory[664]=8'b11111111;
memory[665]=8'b11111111;
memory[666]=8'b11111111;
memory[667]=8'b11111111;
memory[668]=8'b11111111;
memory[669]=8'b11111111;
memory[670]=8'b10000111;
memory[671]=8'b11111111;
memory[672]=8'b11111111;
memory[673]=8'b11111111;
memory[674]=8'b11111111;
memory[675]=8'b11111111;
memory[676]=8'b11111111;
memory[677]=8'b11111111;
memory[678]=8'b11111111;
memory[679]=8'b11111111;
memory[680]=8'b11111111;
memory[681]=8'b11111111;
memory[682]=8'b11111111;
memory[683]=8'b11111111;
memory[684]=8'b11111111;
memory[685]=8'b11111111;
memory[686]=8'b11111111;
memory[687]=8'b11111111;
memory[688]=8'b11111111;
memory[689]=8'b11111111;
memory[690]=8'b11111111;
memory[691]=8'b11111111;
memory[692]=8'b11111111;
memory[693]=8'b11111111;
memory[694]=8'b11111111;
memory[695]=8'b11111111;
memory[696]=8'b11111111;
memory[697]=8'b11111111;
memory[698]=8'b11111111;
memory[699]=8'b11111111;
memory[700]=8'b11110000;
memory[701]=8'b00000000;
memory[702]=8'b00000000;
memory[703]=8'b00000111;
memory[704]=8'b11111111;
memory[705]=8'b11111111;
memory[706]=8'b11111111;
memory[707]=8'b11111111;
memory[708]=8'b11111110;
memory[709]=8'b01111111;
memory[710]=8'b10000011;
memory[711]=8'b11100000;
memory[712]=8'b00011111;
memory[713]=8'b11111111;
memory[714]=8'b11111111;
memory[715]=8'b11111111;
memory[716]=8'b11111111;
memory[717]=8'b11111111;
memory[718]=8'b11111111;
memory[719]=8'b11111111;
memory[720]=8'b11111111;
memory[721]=8'b11111111;
memory[722]=8'b11111111;
memory[723]=8'b11111111;
memory[724]=8'b11111111;
memory[725]=8'b11111111;
memory[726]=8'b11111111;
memory[727]=8'b11111111;
memory[728]=8'b11111111;
memory[729]=8'b11111111;
memory[730]=8'b11111111;
memory[731]=8'b11111111;
memory[732]=8'b11111111;
memory[733]=8'b11111111;
memory[734]=8'b11111111;
memory[735]=8'b11111111;
memory[736]=8'b11111111;
memory[737]=8'b11111111;
memory[738]=8'b11111111;
memory[739]=8'b11111111;
memory[740]=8'b11110000;
memory[741]=8'b00000000;
memory[742]=8'b00000000;
memory[743]=8'b00000111;
memory[744]=8'b11111111;
memory[745]=8'b11111111;
memory[746]=8'b11111111;
memory[747]=8'b11111111;
memory[748]=8'b11111000;
memory[749]=8'b00001111;
memory[750]=8'b10000111;
memory[751]=8'b10000000;
memory[752]=8'b11111111;
memory[753]=8'b11111111;
memory[754]=8'b11111111;
memory[755]=8'b11111111;
memory[756]=8'b11111111;
memory[757]=8'b11111111;
memory[758]=8'b11111111;
memory[759]=8'b11111111;
memory[760]=8'b11111111;
memory[761]=8'b11111111;
memory[762]=8'b11111111;
memory[763]=8'b11111111;
memory[764]=8'b11111111;
memory[765]=8'b11111111;
memory[766]=8'b11111111;
memory[767]=8'b11111111;
memory[768]=8'b11111111;
memory[769]=8'b11111111;
memory[770]=8'b11111111;
memory[771]=8'b11111111;
memory[772]=8'b11111111;
memory[773]=8'b11111111;
memory[774]=8'b11111111;
memory[775]=8'b11111111;
memory[776]=8'b11111111;
memory[777]=8'b11111111;
memory[778]=8'b11111111;
memory[779]=8'b11111111;
memory[780]=8'b11110000;
memory[781]=8'b00000000;
memory[782]=8'b00000000;
memory[783]=8'b00000111;
memory[784]=8'b11111111;
memory[785]=8'b11111111;
memory[786]=8'b11111111;
memory[787]=8'b11111111;
memory[788]=8'b11111100;
memory[789]=8'b00000011;
memory[790]=8'b10000111;
memory[791]=8'b00000001;
memory[792]=8'b11111111;
memory[793]=8'b11111111;
memory[794]=8'b11111111;
memory[795]=8'b11111111;
memory[796]=8'b11111111;
memory[797]=8'b11111111;
memory[798]=8'b11111111;
memory[799]=8'b11111111;
memory[800]=8'b11111111;
memory[801]=8'b11111111;
memory[802]=8'b11111111;
memory[803]=8'b11111111;
memory[804]=8'b11111111;
memory[805]=8'b11111111;
memory[806]=8'b11111111;
memory[807]=8'b11111111;
memory[808]=8'b11111111;
memory[809]=8'b11111111;
memory[810]=8'b11111111;
memory[811]=8'b11111111;
memory[812]=8'b11111111;
memory[813]=8'b11111111;
memory[814]=8'b11111111;
memory[815]=8'b11111111;
memory[816]=8'b11111111;
memory[817]=8'b11111111;
memory[818]=8'b11111111;
memory[819]=8'b11111111;
memory[820]=8'b11111000;
memory[821]=8'b00000000;
memory[822]=8'b00000000;
memory[823]=8'b00001111;
memory[824]=8'b11111111;
memory[825]=8'b11111111;
memory[826]=8'b11111111;
memory[827]=8'b11111111;
memory[828]=8'b11111111;
memory[829]=8'b00000000;
memory[830]=8'b11000100;
memory[831]=8'b00000000;
memory[832]=8'b00001111;
memory[833]=8'b11111111;
memory[834]=8'b11111111;
memory[835]=8'b11111111;
memory[836]=8'b11111111;
memory[837]=8'b11111111;
memory[838]=8'b11111111;
memory[839]=8'b11111111;
memory[840]=8'b11111111;
memory[841]=8'b11111111;
memory[842]=8'b11111111;
memory[843]=8'b11111111;
memory[844]=8'b11111111;
memory[845]=8'b11111111;
memory[846]=8'b11111111;
memory[847]=8'b11111111;
memory[848]=8'b11111111;
memory[849]=8'b11111111;
memory[850]=8'b11111111;
memory[851]=8'b11111111;
memory[852]=8'b11111111;
memory[853]=8'b11111111;
memory[854]=8'b11111111;
memory[855]=8'b11111111;
memory[856]=8'b11111111;
memory[857]=8'b11111111;
memory[858]=8'b11111111;
memory[859]=8'b11111111;
memory[860]=8'b11111000;
memory[861]=8'b00000000;
memory[862]=8'b00000000;
memory[863]=8'b00011111;
memory[864]=8'b11111111;
memory[865]=8'b11111111;
memory[866]=8'b11111111;
memory[867]=8'b11111111;
memory[868]=8'b11111111;
memory[869]=8'b11111100;
memory[870]=8'b01100100;
memory[871]=8'b00000001;
memory[872]=8'b11111111;
memory[873]=8'b11111111;
memory[874]=8'b11111111;
memory[875]=8'b11111111;
memory[876]=8'b11111111;
memory[877]=8'b11111111;
memory[878]=8'b11111111;
memory[879]=8'b11111111;
memory[880]=8'b11111111;
memory[881]=8'b11111111;
memory[882]=8'b11111111;
memory[883]=8'b11111111;
memory[884]=8'b11111111;
memory[885]=8'b11111111;
memory[886]=8'b11111111;
memory[887]=8'b11111111;
memory[888]=8'b11111111;
memory[889]=8'b11111111;
memory[890]=8'b11111111;
memory[891]=8'b11111111;
memory[892]=8'b11111111;
memory[893]=8'b11111111;
memory[894]=8'b11111111;
memory[895]=8'b11111111;
memory[896]=8'b11111111;
memory[897]=8'b11111111;
memory[898]=8'b11111111;
memory[899]=8'b11111111;
memory[900]=8'b11111100;
memory[901]=8'b00000000;
memory[902]=8'b00000000;
memory[903]=8'b00111111;
memory[904]=8'b11111111;
memory[905]=8'b11111111;
memory[906]=8'b11111111;
memory[907]=8'b11111111;
memory[908]=8'b11110000;
memory[909]=8'b00011111;
memory[910]=8'b00100100;
memory[911]=8'b00011111;
memory[912]=8'b11111111;
memory[913]=8'b11111111;
memory[914]=8'b11111111;
memory[915]=8'b11111111;
memory[916]=8'b11111111;
memory[917]=8'b11111111;
memory[918]=8'b11111111;
memory[919]=8'b11111111;
memory[920]=8'b11111111;
memory[921]=8'b11111111;
memory[922]=8'b11111111;
memory[923]=8'b11111111;
memory[924]=8'b11111111;
memory[925]=8'b11111111;
memory[926]=8'b11111111;
memory[927]=8'b11111111;
memory[928]=8'b11111111;
memory[929]=8'b11111111;
memory[930]=8'b11111111;
memory[931]=8'b11111111;
memory[932]=8'b11111111;
memory[933]=8'b11111111;
memory[934]=8'b11111111;
memory[935]=8'b11111111;
memory[936]=8'b11111111;
memory[937]=8'b11111111;
memory[938]=8'b11111111;
memory[939]=8'b11111111;
memory[940]=8'b11111111;
memory[941]=8'b00000000;
memory[942]=8'b00000000;
memory[943]=8'b01111111;
memory[944]=8'b11111111;
memory[945]=8'b11111111;
memory[946]=8'b11111111;
memory[947]=8'b11111111;
memory[948]=8'b10000000;
memory[949]=8'b00000000;
memory[950]=8'b11111111;
memory[951]=8'b11110000;
memory[952]=8'b00000111;
memory[953]=8'b11111111;
memory[954]=8'b11111111;
memory[955]=8'b11111111;
memory[956]=8'b11111111;
memory[957]=8'b11111111;
memory[958]=8'b11111111;
memory[959]=8'b11111111;
memory[960]=8'b11111111;
memory[961]=8'b11111111;
memory[962]=8'b11111111;
memory[963]=8'b11111111;
memory[964]=8'b11111111;
memory[965]=8'b11111111;
memory[966]=8'b11111111;
memory[967]=8'b11111111;
memory[968]=8'b11111111;
memory[969]=8'b11111111;
memory[970]=8'b11111111;
memory[971]=8'b11111111;
memory[972]=8'b11111111;
memory[973]=8'b11111111;
memory[974]=8'b11111111;
memory[975]=8'b11111111;
memory[976]=8'b11111111;
memory[977]=8'b11111111;
memory[978]=8'b11111111;
memory[979]=8'b11111111;
memory[980]=8'b11111111;
memory[981]=8'b11000000;
memory[982]=8'b00000001;
memory[983]=8'b11111111;
memory[984]=8'b11111111;
memory[985]=8'b11111111;
memory[986]=8'b11111111;
memory[987]=8'b11111110;
memory[988]=8'b00000000;
memory[989]=8'b00001110;
memory[990]=8'b01111111;
memory[991]=8'b10000000;
memory[992]=8'b00000001;
memory[993]=8'b11111111;
memory[994]=8'b11111111;
memory[995]=8'b11111111;
memory[996]=8'b11111111;
memory[997]=8'b11111111;
memory[998]=8'b11111111;
memory[999]=8'b11111111;
memory[1000]=8'b11111111;
memory[1001]=8'b11111111;
memory[1002]=8'b11111111;
memory[1003]=8'b11111111;
memory[1004]=8'b11111111;
memory[1005]=8'b11111111;
memory[1006]=8'b11111111;
memory[1007]=8'b11111111;
memory[1008]=8'b11111111;
memory[1009]=8'b11111111;
memory[1010]=8'b11111111;
memory[1011]=8'b11111111;
memory[1012]=8'b11111111;
memory[1013]=8'b11111111;
memory[1014]=8'b11111111;
memory[1015]=8'b11111111;
memory[1016]=8'b11111111;
memory[1017]=8'b11111111;
memory[1018]=8'b11111111;
memory[1019]=8'b11111111;
memory[1020]=8'b11111111;
memory[1021]=8'b11111100;
memory[1022]=8'b00011111;
memory[1023]=8'b11111111;
memory[1024]=8'b11111111;
memory[1025]=8'b11111001;
memory[1026]=8'b11111111;
memory[1027]=8'b11111111;
memory[1028]=8'b11111111;
memory[1029]=8'b00000000;
memory[1030]=8'b00011111;
memory[1031]=8'b10110001;
memory[1032]=8'b11111111;
memory[1033]=8'b11111111;
memory[1034]=8'b11111111;
memory[1035]=8'b11111111;
memory[1036]=8'b11111111;
memory[1037]=8'b11111111;
memory[1038]=8'b11111111;
memory[1039]=8'b11111111;
memory[1040]=8'b11111111;
memory[1041]=8'b11111111;
memory[1042]=8'b11111111;
memory[1043]=8'b11111111;
memory[1044]=8'b11111111;
memory[1045]=8'b11111111;
memory[1046]=8'b11111111;
memory[1047]=8'b11111111;
memory[1048]=8'b11111111;
memory[1049]=8'b11111111;
memory[1050]=8'b11111111;
memory[1051]=8'b11111111;
memory[1052]=8'b11111111;
memory[1053]=8'b11111111;
memory[1054]=8'b11111111;
memory[1055]=8'b11111111;
memory[1056]=8'b11111111;
memory[1057]=8'b11111111;
memory[1058]=8'b11111111;
memory[1059]=8'b11111111;
memory[1060]=8'b11111111;
memory[1061]=8'b11111111;
memory[1062]=8'b11111111;
memory[1063]=8'b11111111;
memory[1064]=8'b11111111;
memory[1065]=8'b10000011;
memory[1066]=8'b11111111;
memory[1067]=8'b11111111;
memory[1068]=8'b11111000;
memory[1069]=8'b00000000;
memory[1070]=8'b00000000;
memory[1071]=8'b00000001;
memory[1072]=8'b11111111;
memory[1073]=8'b11111111;
memory[1074]=8'b11111111;
memory[1075]=8'b11111111;
memory[1076]=8'b11111111;
memory[1077]=8'b11111111;
memory[1078]=8'b11111111;
memory[1079]=8'b11111111;
memory[1080]=8'b11111111;
memory[1081]=8'b11111111;
memory[1082]=8'b11111111;
memory[1083]=8'b11111111;
memory[1084]=8'b11111111;
memory[1085]=8'b11111111;
memory[1086]=8'b11111111;
memory[1087]=8'b11111111;
memory[1088]=8'b11111111;
memory[1089]=8'b11111111;
memory[1090]=8'b11111111;
memory[1091]=8'b11111111;
memory[1092]=8'b11111111;
memory[1093]=8'b11111111;
memory[1094]=8'b11111111;
memory[1095]=8'b11111111;
memory[1096]=8'b11111111;
memory[1097]=8'b11111111;
memory[1098]=8'b11111111;
memory[1099]=8'b11111111;
memory[1100]=8'b11111111;
memory[1101]=8'b11111111;
memory[1102]=8'b11111111;
memory[1103]=8'b11111111;
memory[1104]=8'b11111110;
memory[1105]=8'b00000111;
memory[1106]=8'b11111111;
memory[1107]=8'b11111111;
memory[1108]=8'b11100000;
memory[1109]=8'b10000001;
memory[1110]=8'b00000001;
memory[1111]=8'b10000000;
memory[1112]=8'b11111111;
memory[1113]=8'b11111111;
memory[1114]=8'b11111111;
memory[1115]=8'b11111111;
memory[1116]=8'b11111111;
memory[1117]=8'b11111111;
memory[1118]=8'b11111111;
memory[1119]=8'b11111111;
memory[1120]=8'b11111111;
memory[1121]=8'b11111111;
memory[1122]=8'b11111111;
memory[1123]=8'b11111111;
memory[1124]=8'b11111111;
memory[1125]=8'b11111111;
memory[1126]=8'b11111111;
memory[1127]=8'b11111111;
memory[1128]=8'b11111111;
memory[1129]=8'b11111111;
memory[1130]=8'b11111111;
memory[1131]=8'b11111111;
memory[1132]=8'b11111111;
memory[1133]=8'b11111111;
memory[1134]=8'b11111111;
memory[1135]=8'b11111111;
memory[1136]=8'b11111111;
memory[1137]=8'b11111111;
memory[1138]=8'b11111111;
memory[1139]=8'b11111111;
memory[1140]=8'b11111111;
memory[1141]=8'b11111111;
memory[1142]=8'b11111111;
memory[1143]=8'b11111111;
memory[1144]=8'b11111100;
memory[1145]=8'b00011110;
memory[1146]=8'b00000000;
memory[1147]=8'b11111111;
memory[1148]=8'b10001111;
memory[1149]=8'b11000000;
memory[1150]=8'b00000001;
memory[1151]=8'b10000000;
memory[1152]=8'b00011111;
memory[1153]=8'b11111111;
memory[1154]=8'b11111111;
memory[1155]=8'b11111111;
memory[1156]=8'b11111111;
memory[1157]=8'b11111111;
memory[1158]=8'b11111111;
memory[1159]=8'b11111111;
memory[1160]=8'b11111111;
memory[1161]=8'b11111111;
memory[1162]=8'b11111111;
memory[1163]=8'b11111111;
memory[1164]=8'b11111111;
memory[1165]=8'b11111111;
memory[1166]=8'b11111111;
memory[1167]=8'b11111111;
memory[1168]=8'b11111111;
memory[1169]=8'b11111111;
memory[1170]=8'b11111111;
memory[1171]=8'b11111111;
memory[1172]=8'b11111111;
memory[1173]=8'b11111111;
memory[1174]=8'b11111111;
memory[1175]=8'b11111111;
memory[1176]=8'b11111111;
memory[1177]=8'b11111111;
memory[1178]=8'b11111111;
memory[1179]=8'b11111111;
memory[1180]=8'b11111111;
memory[1181]=8'b11111111;
memory[1182]=8'b11111111;
memory[1183]=8'b11111111;
memory[1184]=8'b11111100;
memory[1185]=8'b00011000;
memory[1186]=8'b00000000;
memory[1187]=8'b00111111;
memory[1188]=8'b11111111;
memory[1189]=8'b10000001;
memory[1190]=8'b10000000;
memory[1191]=8'b11000000;
memory[1192]=8'b00001111;
memory[1193]=8'b11111111;
memory[1194]=8'b11111111;
memory[1195]=8'b11111111;
memory[1196]=8'b11111111;
memory[1197]=8'b11111111;
memory[1198]=8'b11111111;
memory[1199]=8'b11111111;
memory[1200]=8'b11111111;
memory[1201]=8'b11111111;
memory[1202]=8'b11111111;
memory[1203]=8'b11111111;
memory[1204]=8'b11111111;
memory[1205]=8'b11111111;
memory[1206]=8'b11111111;
memory[1207]=8'b11111111;
memory[1208]=8'b11111111;
memory[1209]=8'b11111111;
memory[1210]=8'b11111111;
memory[1211]=8'b11111111;
memory[1212]=8'b11111111;
memory[1213]=8'b11111111;
memory[1214]=8'b11111111;
memory[1215]=8'b11111111;
memory[1216]=8'b11111111;
memory[1217]=8'b11111111;
memory[1218]=8'b11111111;
memory[1219]=8'b11111111;
memory[1220]=8'b11111111;
memory[1221]=8'b11111111;
memory[1222]=8'b11111111;
memory[1223]=8'b11111111;
memory[1224]=8'b11111110;
memory[1225]=8'b00110000;
memory[1226]=8'b01111111;
memory[1227]=8'b00001111;
memory[1228]=8'b11111110;
memory[1229]=8'b00000011;
memory[1230]=8'b10000000;
memory[1231]=8'b11000000;
memory[1232]=8'b00000111;
memory[1233]=8'b11111111;
memory[1234]=8'b11111111;
memory[1235]=8'b11111111;
memory[1236]=8'b11111111;
memory[1237]=8'b11111111;
memory[1238]=8'b11111111;
memory[1239]=8'b11111111;
memory[1240]=8'b11111111;
memory[1241]=8'b11111111;
memory[1242]=8'b11111111;
memory[1243]=8'b11111111;
memory[1244]=8'b11111111;
memory[1245]=8'b11111111;
memory[1246]=8'b11111111;
memory[1247]=8'b11111111;
memory[1248]=8'b11111111;
memory[1249]=8'b11111111;
memory[1250]=8'b11111111;
memory[1251]=8'b11111111;
memory[1252]=8'b11111111;
memory[1253]=8'b11111111;
memory[1254]=8'b11111111;
memory[1255]=8'b11111111;
memory[1256]=8'b11111111;
memory[1257]=8'b11111111;
memory[1258]=8'b11111111;
memory[1259]=8'b11111111;
memory[1260]=8'b11111111;
memory[1261]=8'b11111111;
memory[1262]=8'b11111111;
memory[1263]=8'b11111110;
memory[1264]=8'b00000111;
memory[1265]=8'b00110111;
memory[1266]=8'b11001100;
memory[1267]=8'b01111111;
memory[1268]=8'b11111110;
memory[1269]=8'b00000110;
memory[1270]=8'b01110000;
memory[1271]=8'b11000001;
memory[1272]=8'b00000111;
memory[1273]=8'b11111111;
memory[1274]=8'b11111111;
memory[1275]=8'b11111111;
memory[1276]=8'b11111111;
memory[1277]=8'b11111111;
memory[1278]=8'b11111111;
memory[1279]=8'b11111111;
memory[1280]=8'b11111111;
memory[1281]=8'b11111111;
memory[1282]=8'b11111111;
memory[1283]=8'b11111111;
memory[1284]=8'b11111111;
memory[1285]=8'b11111111;
memory[1286]=8'b11111111;
memory[1287]=8'b11111111;
memory[1288]=8'b11111111;
memory[1289]=8'b11111111;
memory[1290]=8'b11111111;
memory[1291]=8'b11111111;
memory[1292]=8'b11111111;
memory[1293]=8'b11111111;
memory[1294]=8'b11111111;
memory[1295]=8'b11111111;
memory[1296]=8'b11111111;
memory[1297]=8'b11111111;
memory[1298]=8'b11111111;
memory[1299]=8'b11111111;
memory[1300]=8'b11111111;
memory[1301]=8'b11111111;
memory[1302]=8'b11111111;
memory[1303]=8'b11110000;
memory[1304]=8'b00000001;
memory[1305]=8'b10110000;
memory[1306]=8'b00000000;
memory[1307]=8'b00011111;
memory[1308]=8'b11111110;
memory[1309]=8'b00111100;
memory[1310]=8'b01110000;
memory[1311]=8'b01000001;
memory[1312]=8'b11000011;
memory[1313]=8'b11111111;
memory[1314]=8'b11111111;
memory[1315]=8'b11111111;
memory[1316]=8'b11111111;
memory[1317]=8'b11111111;
memory[1318]=8'b11111111;
memory[1319]=8'b11111111;
memory[1320]=8'b11111111;
memory[1321]=8'b11111111;
memory[1322]=8'b11111111;
memory[1323]=8'b11111111;
memory[1324]=8'b11111111;
memory[1325]=8'b11111111;
memory[1326]=8'b11111111;
memory[1327]=8'b11111111;
memory[1328]=8'b11111111;
memory[1329]=8'b11111111;
memory[1330]=8'b11111111;
memory[1331]=8'b11111111;
memory[1332]=8'b11111111;
memory[1333]=8'b11111111;
memory[1334]=8'b11111111;
memory[1335]=8'b11111111;
memory[1336]=8'b11111111;
memory[1337]=8'b11111111;
memory[1338]=8'b11111111;
memory[1339]=8'b11111111;
memory[1340]=8'b11111111;
memory[1341]=8'b11111111;
memory[1342]=8'b11111111;
memory[1343]=8'b11100000;
memory[1344]=8'b00011111;
memory[1345]=8'b11111000;
memory[1346]=8'b00000000;
memory[1347]=8'b00000111;
memory[1348]=8'b11111111;
memory[1349]=8'b11111100;
memory[1350]=8'b11111000;
memory[1351]=8'b01100000;
memory[1352]=8'b11111001;
memory[1353]=8'b11111111;
memory[1354]=8'b11111111;
memory[1355]=8'b11111111;
memory[1356]=8'b11111111;
memory[1357]=8'b11111111;
memory[1358]=8'b11111111;
memory[1359]=8'b11111111;
memory[1360]=8'b11111111;
memory[1361]=8'b11111111;
memory[1362]=8'b11111111;
memory[1363]=8'b11111111;
memory[1364]=8'b11111111;
memory[1365]=8'b11111111;
memory[1366]=8'b11111111;
memory[1367]=8'b11111111;
memory[1368]=8'b11111111;
memory[1369]=8'b11111111;
memory[1370]=8'b11111111;
memory[1371]=8'b11111111;
memory[1372]=8'b11111111;
memory[1373]=8'b11111111;
memory[1374]=8'b11111111;
memory[1375]=8'b11111111;
memory[1376]=8'b11111111;
memory[1377]=8'b11111111;
memory[1378]=8'b11111111;
memory[1379]=8'b11111111;
memory[1380]=8'b11111111;
memory[1381]=8'b11111111;
memory[1382]=8'b11111111;
memory[1383]=8'b11000000;
memory[1384]=8'b11111111;
memory[1385]=8'b11111111;
memory[1386]=8'b10000000;
memory[1387]=8'b00000011;
memory[1388]=8'b11111111;
memory[1389]=8'b11111001;
memory[1390]=8'b11111100;
memory[1391]=8'b01110000;
memory[1392]=8'b11111111;
memory[1393]=8'b11111111;
memory[1394]=8'b11111111;
memory[1395]=8'b11111111;
memory[1396]=8'b11111111;
memory[1397]=8'b11111111;
memory[1398]=8'b11111111;
memory[1399]=8'b11111111;
memory[1400]=8'b11111111;
memory[1401]=8'b11111111;
memory[1402]=8'b11111111;
memory[1403]=8'b11111111;
memory[1404]=8'b11111111;
memory[1405]=8'b11111111;
memory[1406]=8'b11111111;
memory[1407]=8'b11111111;
memory[1408]=8'b11111111;
memory[1409]=8'b11111111;
memory[1410]=8'b11111111;
memory[1411]=8'b11111111;
memory[1412]=8'b11111111;
memory[1413]=8'b11111111;
memory[1414]=8'b11111111;
memory[1415]=8'b11111111;
memory[1416]=8'b11111111;
memory[1417]=8'b11111111;
memory[1418]=8'b11111111;
memory[1419]=8'b11111111;
memory[1420]=8'b11111111;
memory[1421]=8'b11111111;
memory[1422]=8'b11111111;
memory[1423]=8'b10000111;
memory[1424]=8'b11000001;
memory[1425]=8'b11000000;
memory[1426]=8'b01100000;
memory[1427]=8'b00000001;
memory[1428]=8'b11111111;
memory[1429]=8'b11110001;
memory[1430]=8'b11111100;
memory[1431]=8'b01111000;
memory[1432]=8'b11111111;
memory[1433]=8'b11111111;
memory[1434]=8'b11111111;
memory[1435]=8'b11111111;
memory[1436]=8'b11111111;
memory[1437]=8'b11111111;
memory[1438]=8'b11111111;
memory[1439]=8'b11111111;
memory[1440]=8'b11111111;
memory[1441]=8'b11111111;
memory[1442]=8'b11111111;
memory[1443]=8'b11111111;
memory[1444]=8'b11111111;
memory[1445]=8'b11111111;
memory[1446]=8'b11111111;
memory[1447]=8'b11111111;
memory[1448]=8'b11111111;
memory[1449]=8'b11111111;
memory[1450]=8'b11111111;
memory[1451]=8'b11111111;
memory[1452]=8'b11111111;
memory[1453]=8'b11111111;
memory[1454]=8'b11111111;
memory[1455]=8'b11111111;
memory[1456]=8'b11111111;
memory[1457]=8'b11111111;
memory[1458]=8'b11100000;
memory[1459]=8'b00000000;
memory[1460]=8'b11111111;
memory[1461]=8'b11111111;
memory[1462]=8'b11111111;
memory[1463]=8'b00000110;
memory[1464]=8'b00000011;
memory[1465]=8'b11000000;
memory[1466]=8'b00111000;
memory[1467]=8'b00111100;
memory[1468]=8'b11111111;
memory[1469]=8'b11110011;
memory[1470]=8'b11111100;
memory[1471]=8'b01111110;
memory[1472]=8'b11111111;
memory[1473]=8'b11111111;
memory[1474]=8'b11111111;
memory[1475]=8'b11111111;
memory[1476]=8'b11111111;
memory[1477]=8'b11111111;
memory[1478]=8'b11111111;
memory[1479]=8'b11111111;
memory[1480]=8'b11111111;
memory[1481]=8'b11111111;
memory[1482]=8'b11111111;
memory[1483]=8'b11111111;
memory[1484]=8'b11111111;
memory[1485]=8'b11111111;
memory[1486]=8'b11111111;
memory[1487]=8'b11111111;
memory[1488]=8'b11111111;
memory[1489]=8'b11111111;
memory[1490]=8'b11111111;
memory[1491]=8'b11111111;
memory[1492]=8'b11111111;
memory[1493]=8'b11111111;
memory[1494]=8'b11111111;
memory[1495]=8'b11111111;
memory[1496]=8'b11111111;
memory[1497]=8'b11111110;
memory[1498]=8'b00000000;
memory[1499]=8'b00000000;
memory[1500]=8'b00011111;
memory[1501]=8'b11111111;
memory[1502]=8'b11111111;
memory[1503]=8'b00011100;
memory[1504]=8'b00001100;
memory[1505]=8'b00100000;
memory[1506]=8'b00011100;
memory[1507]=8'b00011111;
memory[1508]=8'b11111111;
memory[1509]=8'b11100111;
memory[1510]=8'b11111100;
memory[1511]=8'b01111111;
memory[1512]=8'b11111111;
memory[1513]=8'b11111111;
memory[1514]=8'b11111111;
memory[1515]=8'b11111111;
memory[1516]=8'b11111111;
memory[1517]=8'b11111111;
memory[1518]=8'b11111111;
memory[1519]=8'b11111111;
memory[1520]=8'b11111111;
memory[1521]=8'b11111111;
memory[1522]=8'b11111111;
memory[1523]=8'b11111111;
memory[1524]=8'b11111111;
memory[1525]=8'b11111111;
memory[1526]=8'b11111111;
memory[1527]=8'b11111111;
memory[1528]=8'b11111111;
memory[1529]=8'b11111111;
memory[1530]=8'b11111111;
memory[1531]=8'b11111111;
memory[1532]=8'b11111111;
memory[1533]=8'b11111111;
memory[1534]=8'b11111111;
memory[1535]=8'b11111111;
memory[1536]=8'b11111111;
memory[1537]=8'b11111100;
memory[1538]=8'b00000000;
memory[1539]=8'b00000000;
memory[1540]=8'b00001111;
memory[1541]=8'b11111111;
memory[1542]=8'b11111111;
memory[1543]=8'b00111000;
memory[1544]=8'b00001000;
memory[1545]=8'b00110000;
memory[1546]=8'b00011100;
memory[1547]=8'b00000111;
memory[1548]=8'b11111111;
memory[1549]=8'b11000111;
memory[1550]=8'b11111100;
memory[1551]=8'b11111111;
memory[1552]=8'b11111111;
memory[1553]=8'b11111111;
memory[1554]=8'b11111111;
memory[1555]=8'b11111111;
memory[1556]=8'b11111111;
memory[1557]=8'b11111111;
memory[1558]=8'b11111111;
memory[1559]=8'b11111111;
memory[1560]=8'b11111111;
memory[1561]=8'b11111111;
memory[1562]=8'b11111111;
memory[1563]=8'b11111111;
memory[1564]=8'b11111111;
memory[1565]=8'b11111111;
memory[1566]=8'b11111111;
memory[1567]=8'b11111111;
memory[1568]=8'b11111111;
memory[1569]=8'b11111111;
memory[1570]=8'b11111111;
memory[1571]=8'b11111111;
memory[1572]=8'b11111111;
memory[1573]=8'b11111111;
memory[1574]=8'b11111111;
memory[1575]=8'b11111111;
memory[1576]=8'b11111111;
memory[1577]=8'b11111000;
memory[1578]=8'b00000000;
memory[1579]=8'b00111110;
memory[1580]=8'b00001111;
memory[1581]=8'b11111111;
memory[1582]=8'b11111110;
memory[1583]=8'b01111000;
memory[1584]=8'b00000000;
memory[1585]=8'b00011000;
memory[1586]=8'b00000001;
memory[1587]=8'b00000011;
memory[1588]=8'b11111111;
memory[1589]=8'b11001111;
memory[1590]=8'b11111111;
memory[1591]=8'b11111111;
memory[1592]=8'b11111111;
memory[1593]=8'b11111111;
memory[1594]=8'b11111111;
memory[1595]=8'b11111111;
memory[1596]=8'b11111111;
memory[1597]=8'b11111111;
memory[1598]=8'b11111111;
memory[1599]=8'b11111111;
memory[1600]=8'b11111111;
memory[1601]=8'b11111111;
memory[1602]=8'b11111111;
memory[1603]=8'b11111111;
memory[1604]=8'b11111111;
memory[1605]=8'b11111111;
memory[1606]=8'b11111111;
memory[1607]=8'b11111111;
memory[1608]=8'b11111111;
memory[1609]=8'b11111111;
memory[1610]=8'b11111111;
memory[1611]=8'b11111111;
memory[1612]=8'b11111111;
memory[1613]=8'b11111111;
memory[1614]=8'b11111111;
memory[1615]=8'b11111111;
memory[1616]=8'b11111111;
memory[1617]=8'b11110000;
memory[1618]=8'b00000000;
memory[1619]=8'b01110111;
memory[1620]=8'b11111111;
memory[1621]=8'b11111111;
memory[1622]=8'b11111111;
memory[1623]=8'b11110000;
memory[1624]=8'b00000000;
memory[1625]=8'b00011000;
memory[1626]=8'b00000001;
memory[1627]=8'b11000001;
memory[1628]=8'b11111111;
memory[1629]=8'b10001111;
memory[1630]=8'b11111111;
memory[1631]=8'b11111111;
memory[1632]=8'b11111111;
memory[1633]=8'b11111111;
memory[1634]=8'b11111111;
memory[1635]=8'b11111111;
memory[1636]=8'b11111111;
memory[1637]=8'b11111111;
memory[1638]=8'b11111111;
memory[1639]=8'b11111111;
memory[1640]=8'b11111111;
memory[1641]=8'b11111111;
memory[1642]=8'b11111111;
memory[1643]=8'b11111111;
memory[1644]=8'b11111111;
memory[1645]=8'b11111111;
memory[1646]=8'b11111111;
memory[1647]=8'b11111111;
memory[1648]=8'b11111111;
memory[1649]=8'b11111111;
memory[1650]=8'b11111111;
memory[1651]=8'b11111111;
memory[1652]=8'b11111111;
memory[1653]=8'b11111111;
memory[1654]=8'b11111111;
memory[1655]=8'b11111111;
memory[1656]=8'b11111111;
memory[1657]=8'b11100000;
memory[1658]=8'b00000000;
memory[1659]=8'b01111111;
memory[1660]=8'b11111111;
memory[1661]=8'b11111111;
memory[1662]=8'b11111111;
memory[1663]=8'b11110000;
memory[1664]=8'b00010000;
memory[1665]=8'b00011100;
memory[1666]=8'b00001100;
memory[1667]=8'b11111001;
memory[1668]=8'b11111111;
memory[1669]=8'b00011111;
memory[1670]=8'b11111111;
memory[1671]=8'b11111111;
memory[1672]=8'b11111111;
memory[1673]=8'b11111111;
memory[1674]=8'b11111111;
memory[1675]=8'b11111111;
memory[1676]=8'b11111111;
memory[1677]=8'b11111111;
memory[1678]=8'b11111111;
memory[1679]=8'b11111111;
memory[1680]=8'b11111111;
memory[1681]=8'b11111111;
memory[1682]=8'b11111111;
memory[1683]=8'b11111111;
memory[1684]=8'b11111111;
memory[1685]=8'b11111111;
memory[1686]=8'b11111111;
memory[1687]=8'b11111111;
memory[1688]=8'b11111111;
memory[1689]=8'b11111111;
memory[1690]=8'b11111111;
memory[1691]=8'b11111111;
memory[1692]=8'b11111111;
memory[1693]=8'b11111111;
memory[1694]=8'b11111111;
memory[1695]=8'b11111111;
memory[1696]=8'b11111111;
memory[1697]=8'b11000000;
memory[1698]=8'b00000000;
memory[1699]=8'b00111111;
memory[1700]=8'b11111111;
memory[1701]=8'b11111111;
memory[1702]=8'b11111111;
memory[1703]=8'b11110000;
memory[1704]=8'b01100000;
memory[1705]=8'b00011110;
memory[1706]=8'b00011110;
memory[1707]=8'b01111111;
memory[1708]=8'b11111111;
memory[1709]=8'b00111111;
memory[1710]=8'b11111111;
memory[1711]=8'b11111111;
memory[1712]=8'b11111111;
memory[1713]=8'b11111111;
memory[1714]=8'b11111111;
memory[1715]=8'b11111111;
memory[1716]=8'b11111111;
memory[1717]=8'b11111111;
memory[1718]=8'b11111111;
memory[1719]=8'b11111111;
memory[1720]=8'b11111111;
memory[1721]=8'b11111111;
memory[1722]=8'b11111111;
memory[1723]=8'b11111111;
memory[1724]=8'b11111111;
memory[1725]=8'b11111111;
memory[1726]=8'b11111111;
memory[1727]=8'b11111111;
memory[1728]=8'b11111111;
memory[1729]=8'b11111111;
memory[1730]=8'b11111111;
memory[1731]=8'b11111111;
memory[1732]=8'b11111111;
memory[1733]=8'b11111111;
memory[1734]=8'b11111111;
memory[1735]=8'b11111111;
memory[1736]=8'b11111111;
memory[1737]=8'b11000000;
memory[1738]=8'b00000000;
memory[1739]=8'b00000111;
memory[1740]=8'b11111111;
memory[1741]=8'b11111111;
memory[1742]=8'b11111111;
memory[1743]=8'b11111000;
memory[1744]=8'b01100000;
memory[1745]=8'b00001111;
memory[1746]=8'b00011110;
memory[1747]=8'b00111111;
memory[1748]=8'b11111110;
memory[1749]=8'b00111111;
memory[1750]=8'b11111111;
memory[1751]=8'b11111111;
memory[1752]=8'b11111111;
memory[1753]=8'b11111111;
memory[1754]=8'b11111111;
memory[1755]=8'b11111111;
memory[1756]=8'b11111111;
memory[1757]=8'b11111111;
memory[1758]=8'b11111111;
memory[1759]=8'b11111111;
memory[1760]=8'b11111111;
memory[1761]=8'b11111111;
memory[1762]=8'b11111111;
memory[1763]=8'b11111111;
memory[1764]=8'b11111111;
memory[1765]=8'b11111111;
memory[1766]=8'b11111111;
memory[1767]=8'b11111111;
memory[1768]=8'b11111111;
memory[1769]=8'b11111111;
memory[1770]=8'b11111111;
memory[1771]=8'b11111111;
memory[1772]=8'b11111111;
memory[1773]=8'b11111111;
memory[1774]=8'b11111111;
memory[1775]=8'b11111111;
memory[1776]=8'b11111111;
memory[1777]=8'b10000000;
memory[1778]=8'b00000000;
memory[1779]=8'b00000001;
memory[1780]=8'b11111111;
memory[1781]=8'b11111111;
memory[1782]=8'b11111111;
memory[1783]=8'b11111000;
memory[1784]=8'b01110000;
memory[1785]=8'b00001111;
memory[1786]=8'b10011111;
memory[1787]=8'b00011111;
memory[1788]=8'b11111110;
memory[1789]=8'b00111111;
memory[1790]=8'b11111111;
memory[1791]=8'b11111111;
memory[1792]=8'b11111111;
memory[1793]=8'b11111111;
memory[1794]=8'b11111111;
memory[1795]=8'b11111111;
memory[1796]=8'b11111111;
memory[1797]=8'b11111111;
memory[1798]=8'b11111111;
memory[1799]=8'b11111111;
memory[1800]=8'b11111111;
memory[1801]=8'b11111111;
memory[1802]=8'b11111111;
memory[1803]=8'b11111111;
memory[1804]=8'b11111111;
memory[1805]=8'b11111111;
memory[1806]=8'b11111111;
memory[1807]=8'b11111111;
memory[1808]=8'b11111111;
memory[1809]=8'b11111111;
memory[1810]=8'b11111111;
memory[1811]=8'b11111111;
memory[1812]=8'b11111111;
memory[1813]=8'b11111111;
memory[1814]=8'b11111111;
memory[1815]=8'b11111111;
memory[1816]=8'b11111111;
memory[1817]=8'b10000000;
memory[1818]=8'b00000011;
memory[1819]=8'b11110001;
memory[1820]=8'b11111111;
memory[1821]=8'b11111111;
memory[1822]=8'b11111111;
memory[1823]=8'b11111111;
memory[1824]=8'b11111000;
memory[1825]=8'b00011111;
memory[1826]=8'b11111111;
memory[1827]=8'b10001111;
memory[1828]=8'b11111100;
memory[1829]=8'b01111111;
memory[1830]=8'b11111111;
memory[1831]=8'b11111111;
memory[1832]=8'b11111111;
memory[1833]=8'b11111111;
memory[1834]=8'b11111111;
memory[1835]=8'b11111111;
memory[1836]=8'b11111111;
memory[1837]=8'b11111111;
memory[1838]=8'b11111111;
memory[1839]=8'b11111111;
memory[1840]=8'b11111111;
memory[1841]=8'b11111111;
memory[1842]=8'b11111111;
memory[1843]=8'b11111111;
memory[1844]=8'b11111111;
memory[1845]=8'b11111111;
memory[1846]=8'b11111111;
memory[1847]=8'b11111111;
memory[1848]=8'b11111111;
memory[1849]=8'b11111111;
memory[1850]=8'b11111111;
memory[1851]=8'b11111111;
memory[1852]=8'b11111111;
memory[1853]=8'b11111111;
memory[1854]=8'b11111111;
memory[1855]=8'b11111111;
memory[1856]=8'b11111111;
memory[1857]=8'b10000000;
memory[1858]=8'b00001111;
memory[1859]=8'b11111111;
memory[1860]=8'b11111111;
memory[1861]=8'b11111111;
memory[1862]=8'b11111111;
memory[1863]=8'b11111111;
memory[1864]=8'b11111100;
memory[1865]=8'b00001111;
memory[1866]=8'b11111111;
memory[1867]=8'b11000111;
memory[1868]=8'b11111000;
memory[1869]=8'b01111111;
memory[1870]=8'b11111111;
memory[1871]=8'b11111111;
memory[1872]=8'b11111111;
memory[1873]=8'b11111111;
memory[1874]=8'b11111111;
memory[1875]=8'b11111111;
memory[1876]=8'b11111111;
memory[1877]=8'b11111111;
memory[1878]=8'b11111111;
memory[1879]=8'b11111111;
memory[1880]=8'b11111111;
memory[1881]=8'b11111111;
memory[1882]=8'b11111111;
memory[1883]=8'b11111111;
memory[1884]=8'b11111111;
memory[1885]=8'b11111111;
memory[1886]=8'b11111111;
memory[1887]=8'b11111111;
memory[1888]=8'b11111111;
memory[1889]=8'b11111111;
memory[1890]=8'b11111111;
memory[1891]=8'b11111111;
memory[1892]=8'b11111111;
memory[1893]=8'b11111111;
memory[1894]=8'b11111111;
memory[1895]=8'b11111111;
memory[1896]=8'b11111111;
memory[1897]=8'b10000000;
memory[1898]=8'b00011111;
memory[1899]=8'b11111111;
memory[1900]=8'b11111111;
memory[1901]=8'b11010111;
memory[1902]=8'b11111111;
memory[1903]=8'b11111111;
memory[1904]=8'b11111110;
memory[1905]=8'b00011111;
memory[1906]=8'b11111111;
memory[1907]=8'b11100111;
memory[1908]=8'b11111000;
memory[1909]=8'b01111111;
memory[1910]=8'b11111111;
memory[1911]=8'b11111111;
memory[1912]=8'b11111111;
memory[1913]=8'b11111111;
memory[1914]=8'b11111111;
memory[1915]=8'b11111111;
memory[1916]=8'b11111111;
memory[1917]=8'b11111111;
memory[1918]=8'b11111111;
memory[1919]=8'b11111111;
memory[1920]=8'b11111111;
memory[1921]=8'b11111111;
memory[1922]=8'b11111111;
memory[1923]=8'b11111111;
memory[1924]=8'b11111111;
memory[1925]=8'b11111111;
memory[1926]=8'b11111111;
memory[1927]=8'b11111111;
memory[1928]=8'b11111111;
memory[1929]=8'b11111111;
memory[1930]=8'b11111111;
memory[1931]=8'b11111111;
memory[1932]=8'b11111111;
memory[1933]=8'b11111111;
memory[1934]=8'b11111111;
memory[1935]=8'b11111111;
memory[1936]=8'b11111111;
memory[1937]=8'b00000000;
memory[1938]=8'b00111111;
memory[1939]=8'b11111111;
memory[1940]=8'b11111111;
memory[1941]=8'b10000011;
memory[1942]=8'b11111111;
memory[1943]=8'b11111111;
memory[1944]=8'b11111111;
memory[1945]=8'b00011111;
memory[1946]=8'b11111111;
memory[1947]=8'b11100011;
memory[1948]=8'b11110000;
memory[1949]=8'b01111111;
memory[1950]=8'b11111111;
memory[1951]=8'b11111111;
memory[1952]=8'b11111111;
memory[1953]=8'b11111111;
memory[1954]=8'b11111111;
memory[1955]=8'b11111111;
memory[1956]=8'b11111111;
memory[1957]=8'b11111111;
memory[1958]=8'b11111111;
memory[1959]=8'b11111111;
memory[1960]=8'b11111111;
memory[1961]=8'b11111111;
memory[1962]=8'b11111111;
memory[1963]=8'b11111111;
memory[1964]=8'b11111111;
memory[1965]=8'b11111111;
memory[1966]=8'b11111111;
memory[1967]=8'b11111111;
memory[1968]=8'b11111111;
memory[1969]=8'b11111111;
memory[1970]=8'b11111111;
memory[1971]=8'b11111111;
memory[1972]=8'b11111111;
memory[1973]=8'b11111111;
memory[1974]=8'b11111111;
memory[1975]=8'b11111111;
memory[1976]=8'b11111111;
memory[1977]=8'b00000000;
memory[1978]=8'b00111111;
memory[1979]=8'b11111111;
memory[1980]=8'b11111110;
memory[1981]=8'b00000011;
memory[1982]=8'b11111111;
memory[1983]=8'b11111111;
memory[1984]=8'b11111111;
memory[1985]=8'b10011111;
memory[1986]=8'b11111111;
memory[1987]=8'b11110001;
memory[1988]=8'b11110000;
memory[1989]=8'b11111111;
memory[1990]=8'b11111111;
memory[1991]=8'b11111111;
memory[1992]=8'b11111111;
memory[1993]=8'b11111111;
memory[1994]=8'b11111111;
memory[1995]=8'b11111111;
memory[1996]=8'b11111111;
memory[1997]=8'b11111111;
memory[1998]=8'b11111111;
memory[1999]=8'b11111111;
memory[2000]=8'b11111111;
memory[2001]=8'b11111111;
memory[2002]=8'b11111111;
memory[2003]=8'b11111111;
memory[2004]=8'b11111111;
memory[2005]=8'b11111111;
memory[2006]=8'b11111111;
memory[2007]=8'b11111111;
memory[2008]=8'b11111111;
memory[2009]=8'b11111111;
memory[2010]=8'b11111111;
memory[2011]=8'b11111111;
memory[2012]=8'b11111111;
memory[2013]=8'b11111111;
memory[2014]=8'b11111111;
memory[2015]=8'b11111111;
memory[2016]=8'b11111111;
memory[2017]=8'b10000000;
memory[2018]=8'b00111111;
memory[2019]=8'b11111111;
memory[2020]=8'b11111111;
memory[2021]=8'b00000111;
memory[2022]=8'b11111111;
memory[2023]=8'b11111111;
memory[2024]=8'b11111111;
memory[2025]=8'b11111111;
memory[2026]=8'b11111111;
memory[2027]=8'b11110001;
memory[2028]=8'b11100000;
memory[2029]=8'b11111111;
memory[2030]=8'b11111111;
memory[2031]=8'b11111111;
memory[2032]=8'b11111111;
memory[2033]=8'b11111111;
memory[2034]=8'b11111111;
memory[2035]=8'b11111111;
memory[2036]=8'b11111111;
memory[2037]=8'b11111111;
memory[2038]=8'b11111111;
memory[2039]=8'b11111111;
memory[2040]=8'b11111111;
memory[2041]=8'b11111111;
memory[2042]=8'b11111111;
memory[2043]=8'b11111111;
memory[2044]=8'b11111111;
memory[2045]=8'b11111111;
memory[2046]=8'b11111111;
memory[2047]=8'b11111111;
memory[2048]=8'b11111111;
memory[2049]=8'b11111111;
memory[2050]=8'b11111111;
memory[2051]=8'b11111111;
memory[2052]=8'b11111111;
memory[2053]=8'b11111111;
memory[2054]=8'b11111111;
memory[2055]=8'b11111111;
memory[2056]=8'b11111111;
memory[2057]=8'b10000000;
memory[2058]=8'b00011111;
memory[2059]=8'b11111111;
memory[2060]=8'b11111111;
memory[2061]=8'b00000111;
memory[2062]=8'b11111111;
memory[2063]=8'b11111111;
memory[2064]=8'b11111111;
memory[2065]=8'b11111111;
memory[2066]=8'b11111111;
memory[2067]=8'b11111000;
memory[2068]=8'b11100001;
memory[2069]=8'b11111111;
memory[2070]=8'b11111111;
memory[2071]=8'b11111111;
memory[2072]=8'b11111111;
memory[2073]=8'b11111111;
memory[2074]=8'b11111111;
memory[2075]=8'b11111111;
memory[2076]=8'b11111111;
memory[2077]=8'b11111111;
memory[2078]=8'b11111111;
memory[2079]=8'b11111111;
memory[2080]=8'b11111111;
memory[2081]=8'b11111111;
memory[2082]=8'b11111111;
memory[2083]=8'b11111111;
memory[2084]=8'b11111111;
memory[2085]=8'b11111111;
memory[2086]=8'b11111111;
memory[2087]=8'b11111111;
memory[2088]=8'b11111111;
memory[2089]=8'b11111111;
memory[2090]=8'b11111111;
memory[2091]=8'b11111111;
memory[2092]=8'b11111111;
memory[2093]=8'b11111111;
memory[2094]=8'b11111111;
memory[2095]=8'b11111111;
memory[2096]=8'b11111111;
memory[2097]=8'b10000000;
memory[2098]=8'b00001111;
memory[2099]=8'b11111111;
memory[2100]=8'b11111111;
memory[2101]=8'b10000111;
memory[2102]=8'b11111111;
memory[2103]=8'b11111111;
memory[2104]=8'b11111111;
memory[2105]=8'b11111111;
memory[2106]=8'b11111111;
memory[2107]=8'b11111000;
memory[2108]=8'b11100001;
memory[2109]=8'b11111111;
memory[2110]=8'b11111111;
memory[2111]=8'b11111111;
memory[2112]=8'b11111111;
memory[2113]=8'b11111111;
memory[2114]=8'b11111111;
memory[2115]=8'b11111111;
memory[2116]=8'b11111111;
memory[2117]=8'b11111111;
memory[2118]=8'b11111111;
memory[2119]=8'b11111111;
memory[2120]=8'b11111111;
memory[2121]=8'b11111111;
memory[2122]=8'b11111111;
memory[2123]=8'b11111111;
memory[2124]=8'b11111111;
memory[2125]=8'b11111111;
memory[2126]=8'b11111111;
memory[2127]=8'b11111111;
memory[2128]=8'b11111111;
memory[2129]=8'b11111111;
memory[2130]=8'b11111111;
memory[2131]=8'b11111111;
memory[2132]=8'b11111111;
memory[2133]=8'b11111111;
memory[2134]=8'b11111111;
memory[2135]=8'b11111111;
memory[2136]=8'b11111111;
memory[2137]=8'b11000000;
memory[2138]=8'b00000111;
memory[2139]=8'b11111111;
memory[2140]=8'b11111111;
memory[2141]=8'b11000111;
memory[2142]=8'b11111111;
memory[2143]=8'b11111111;
memory[2144]=8'b11111111;
memory[2145]=8'b11111111;
memory[2146]=8'b11111111;
memory[2147]=8'b11111000;
memory[2148]=8'b01000001;
memory[2149]=8'b11111111;
memory[2150]=8'b11111111;
memory[2151]=8'b11111111;
memory[2152]=8'b11111111;
memory[2153]=8'b11111111;
memory[2154]=8'b11111111;
memory[2155]=8'b11111111;
memory[2156]=8'b11111111;
memory[2157]=8'b11111111;
memory[2158]=8'b11111111;
memory[2159]=8'b11111111;
memory[2160]=8'b11111111;
memory[2161]=8'b11111111;
memory[2162]=8'b11111111;
memory[2163]=8'b11111111;
memory[2164]=8'b11111111;
memory[2165]=8'b11111111;
memory[2166]=8'b11111111;
memory[2167]=8'b11111111;
memory[2168]=8'b11111111;
memory[2169]=8'b11111111;
memory[2170]=8'b11111111;
memory[2171]=8'b11111111;
memory[2172]=8'b11111111;
memory[2173]=8'b11111111;
memory[2174]=8'b11111111;
memory[2175]=8'b11111111;
memory[2176]=8'b11111111;
memory[2177]=8'b11000000;
memory[2178]=8'b00000111;
memory[2179]=8'b11111111;
memory[2180]=8'b11111111;
memory[2181]=8'b11001111;
memory[2182]=8'b11111111;
memory[2183]=8'b11111111;
memory[2184]=8'b11111111;
memory[2185]=8'b11111111;
memory[2186]=8'b11111111;
memory[2187]=8'b11111100;
memory[2188]=8'b00000001;
memory[2189]=8'b11111111;
memory[2190]=8'b11111111;
memory[2191]=8'b11111111;
memory[2192]=8'b11111111;
memory[2193]=8'b11111111;
memory[2194]=8'b11111111;
memory[2195]=8'b11111111;
memory[2196]=8'b11111111;
memory[2197]=8'b11111111;
memory[2198]=8'b11111111;
memory[2199]=8'b11111111;
memory[2200]=8'b11111111;
memory[2201]=8'b11111111;
memory[2202]=8'b11111111;
memory[2203]=8'b11111111;
memory[2204]=8'b11111111;
memory[2205]=8'b11111111;
memory[2206]=8'b11111111;
memory[2207]=8'b11111111;
memory[2208]=8'b11111111;
memory[2209]=8'b11111111;
memory[2210]=8'b11111111;
memory[2211]=8'b11111111;
memory[2212]=8'b11111111;
memory[2213]=8'b11111111;
memory[2214]=8'b11111111;
memory[2215]=8'b11111111;
memory[2216]=8'b11111111;
memory[2217]=8'b11100000;
memory[2218]=8'b00000011;
memory[2219]=8'b11111111;
memory[2220]=8'b11111111;
memory[2221]=8'b11001111;
memory[2222]=8'b11111111;
memory[2223]=8'b11111111;
memory[2224]=8'b11111111;
memory[2225]=8'b11111111;
memory[2226]=8'b11111111;
memory[2227]=8'b11111100;
memory[2228]=8'b00000001;
memory[2229]=8'b11111111;
memory[2230]=8'b11111111;
memory[2231]=8'b11111111;
memory[2232]=8'b11111111;
memory[2233]=8'b11111111;
memory[2234]=8'b11111111;
memory[2235]=8'b11111111;
memory[2236]=8'b11111111;
memory[2237]=8'b11111111;
memory[2238]=8'b11111111;
memory[2239]=8'b11111111;
memory[2240]=8'b11111111;
memory[2241]=8'b11111111;
memory[2242]=8'b11111111;
memory[2243]=8'b11111111;
memory[2244]=8'b11111111;
memory[2245]=8'b11111111;
memory[2246]=8'b11111111;
memory[2247]=8'b11111111;
memory[2248]=8'b11111111;
memory[2249]=8'b11111111;
memory[2250]=8'b11111111;
memory[2251]=8'b11111111;
memory[2252]=8'b11111111;
memory[2253]=8'b11111111;
memory[2254]=8'b11111111;
memory[2255]=8'b11111111;
memory[2256]=8'b11111111;
memory[2257]=8'b11110000;
memory[2258]=8'b00000001;
memory[2259]=8'b11111111;
memory[2260]=8'b11111111;
memory[2261]=8'b11111111;
memory[2262]=8'b11111111;
memory[2263]=8'b11111111;
memory[2264]=8'b11111111;
memory[2265]=8'b11111111;
memory[2266]=8'b11111111;
memory[2267]=8'b11111000;
memory[2268]=8'b00010011;
memory[2269]=8'b11111111;
memory[2270]=8'b11111111;
memory[2271]=8'b11111111;
memory[2272]=8'b11111111;
memory[2273]=8'b11111111;
memory[2274]=8'b11111111;
memory[2275]=8'b11111111;
memory[2276]=8'b11111111;
memory[2277]=8'b11111111;
memory[2278]=8'b11111111;
memory[2279]=8'b11111111;
memory[2280]=8'b11111111;
memory[2281]=8'b11111111;
memory[2282]=8'b11111111;
memory[2283]=8'b11111111;
memory[2284]=8'b11111111;
memory[2285]=8'b11111111;
memory[2286]=8'b11111111;
memory[2287]=8'b11111111;
memory[2288]=8'b11111111;
memory[2289]=8'b11111111;
memory[2290]=8'b11111111;
memory[2291]=8'b11111111;
memory[2292]=8'b11111111;
memory[2293]=8'b11111111;
memory[2294]=8'b11111111;
memory[2295]=8'b11111111;
memory[2296]=8'b11111111;
memory[2297]=8'b11110000;
memory[2298]=8'b00000000;
memory[2299]=8'b11111111;
memory[2300]=8'b11111111;
memory[2301]=8'b11111111;
memory[2302]=8'b11111111;
memory[2303]=8'b11111111;
memory[2304]=8'b11111111;
memory[2305]=8'b11111111;
memory[2306]=8'b11111111;
memory[2307]=8'b00000000;
memory[2308]=8'b00000011;
memory[2309]=8'b11111111;
memory[2310]=8'b11111111;
memory[2311]=8'b11111111;
memory[2312]=8'b11111111;
memory[2313]=8'b11111111;
memory[2314]=8'b11111111;
memory[2315]=8'b11111111;
memory[2316]=8'b11111111;
memory[2317]=8'b11111111;
memory[2318]=8'b11111111;
memory[2319]=8'b11111111;
memory[2320]=8'b11111111;
memory[2321]=8'b11111111;
memory[2322]=8'b11111111;
memory[2323]=8'b11111111;
memory[2324]=8'b11111111;
memory[2325]=8'b11111111;
memory[2326]=8'b11111111;
memory[2327]=8'b11111111;
memory[2328]=8'b11111111;
memory[2329]=8'b11111111;
memory[2330]=8'b11111111;
memory[2331]=8'b11111111;
memory[2332]=8'b11111111;
memory[2333]=8'b11111111;
memory[2334]=8'b11111111;
memory[2335]=8'b11111111;
memory[2336]=8'b11111111;
memory[2337]=8'b11111000;
memory[2338]=8'b00000000;
memory[2339]=8'b01111111;
memory[2340]=8'b11111111;
memory[2341]=8'b11111111;
memory[2342]=8'b11111111;
memory[2343]=8'b11111111;
memory[2344]=8'b11111111;
memory[2345]=8'b11111111;
memory[2346]=8'b11111000;
memory[2347]=8'b00000000;
memory[2348]=8'b00000000;
memory[2349]=8'b01111111;
memory[2350]=8'b11111111;
memory[2351]=8'b11111111;
memory[2352]=8'b11111111;
memory[2353]=8'b11111111;
memory[2354]=8'b11111111;
memory[2355]=8'b11111111;
memory[2356]=8'b11111111;
memory[2357]=8'b11111111;
memory[2358]=8'b11111111;
memory[2359]=8'b11111111;
memory[2360]=8'b11111111;
memory[2361]=8'b11111111;
memory[2362]=8'b11111111;
memory[2363]=8'b11111111;
memory[2364]=8'b11111111;
memory[2365]=8'b11111111;
memory[2366]=8'b11111111;
memory[2367]=8'b11111111;
memory[2368]=8'b11111111;
memory[2369]=8'b11111111;
memory[2370]=8'b11111111;
memory[2371]=8'b11111111;
memory[2372]=8'b11111111;
memory[2373]=8'b11111111;
memory[2374]=8'b11111111;
memory[2375]=8'b11111111;
memory[2376]=8'b11111111;
memory[2377]=8'b11111100;
memory[2378]=8'b00000000;
memory[2379]=8'b00111111;
memory[2380]=8'b11111111;
memory[2381]=8'b11111111;
memory[2382]=8'b11111111;
memory[2383]=8'b11111111;
memory[2384]=8'b11111111;
memory[2385]=8'b11111111;
memory[2386]=8'b11000000;
memory[2387]=8'b00000000;
memory[2388]=8'b00000000;
memory[2389]=8'b00001111;
memory[2390]=8'b11111111;
memory[2391]=8'b11111111;
memory[2392]=8'b11111111;
memory[2393]=8'b11111111;
memory[2394]=8'b11111111;
memory[2395]=8'b11111111;
memory[2396]=8'b11111111;
memory[2397]=8'b11111111;
memory[2398]=8'b11111111;
memory[2399]=8'b11111111;
memory[2400]=8'b11111111;
memory[2401]=8'b11111111;
memory[2402]=8'b11111111;
memory[2403]=8'b11111111;
memory[2404]=8'b11111111;
memory[2405]=8'b11111111;
memory[2406]=8'b11111111;
memory[2407]=8'b11111111;
memory[2408]=8'b10000000;
memory[2409]=8'b00000000;
memory[2410]=8'b00000000;
memory[2411]=8'b00000000;
memory[2412]=8'b00000000;
memory[2413]=8'b00000000;
memory[2414]=8'b00000000;
memory[2415]=8'b00000000;
memory[2416]=8'b00000011;
memory[2417]=8'b11111110;
memory[2418]=8'b00000000;
memory[2419]=8'b00011111;
memory[2420]=8'b11111111;
memory[2421]=8'b11100000;
memory[2422]=8'b00000000;
memory[2423]=8'b00011111;
memory[2424]=8'b11111111;
memory[2425]=8'b11111111;
memory[2426]=8'b00000000;
memory[2427]=8'b00000000;
memory[2428]=8'b00000000;
memory[2429]=8'b00000011;
memory[2430]=8'b11111111;
memory[2431]=8'b11111111;
memory[2432]=8'b11111111;
memory[2433]=8'b11111111;
memory[2434]=8'b11111111;
memory[2435]=8'b11111111;
memory[2436]=8'b11111111;
memory[2437]=8'b11111111;
memory[2438]=8'b11111111;
memory[2439]=8'b11111111;
memory[2440]=8'b11111111;
memory[2441]=8'b11111111;
memory[2442]=8'b11111111;
memory[2443]=8'b11111111;
memory[2444]=8'b11111111;
memory[2445]=8'b11111111;
memory[2446]=8'b11111111;
memory[2447]=8'b11111111;
memory[2448]=8'b11111000;
memory[2449]=8'b00000000;
memory[2450]=8'b00111111;
memory[2451]=8'b11111111;
memory[2452]=8'b00000000;
memory[2453]=8'b00111111;
memory[2454]=8'b11111110;
memory[2455]=8'b00000011;
memory[2456]=8'b11111111;
memory[2457]=8'b11111111;
memory[2458]=8'b00000000;
memory[2459]=8'b00001111;
memory[2460]=8'b11111111;
memory[2461]=8'b11111111;
memory[2462]=8'b11111111;
memory[2463]=8'b11111111;
memory[2464]=8'b11111111;
memory[2465]=8'b11111000;
memory[2466]=8'b00000000;
memory[2467]=8'b00000000;
memory[2468]=8'b00000000;
memory[2469]=8'b00000000;
memory[2470]=8'b11111111;
memory[2471]=8'b11111111;
memory[2472]=8'b11111111;
memory[2473]=8'b11111111;
memory[2474]=8'b11111111;
memory[2475]=8'b11111111;
memory[2476]=8'b11111111;
memory[2477]=8'b11111111;
memory[2478]=8'b11111111;
memory[2479]=8'b11111111;
memory[2480]=8'b11111111;
memory[2481]=8'b11111111;
memory[2482]=8'b11111111;
memory[2483]=8'b11111111;
memory[2484]=8'b11111111;
memory[2485]=8'b11111111;
memory[2486]=8'b11111111;
memory[2487]=8'b11111111;
memory[2488]=8'b11111111;
memory[2489]=8'b11111111;
memory[2490]=8'b11111111;
memory[2491]=8'b11111111;
memory[2492]=8'b11111111;
memory[2493]=8'b11111111;
memory[2494]=8'b11111111;
memory[2495]=8'b11111111;
memory[2496]=8'b11111111;
memory[2497]=8'b11111111;
memory[2498]=8'b10000000;
memory[2499]=8'b00000111;
memory[2500]=8'b11111111;
memory[2501]=8'b11111111;
memory[2502]=8'b11111111;
memory[2503]=8'b11111111;
memory[2504]=8'b11111111;
memory[2505]=8'b10000000;
memory[2506]=8'b00000000;
memory[2507]=8'b00000000;
memory[2508]=8'b00000000;
memory[2509]=8'b00000000;
memory[2510]=8'b00111111;
memory[2511]=8'b11111111;
memory[2512]=8'b11111111;
memory[2513]=8'b11111111;
memory[2514]=8'b11111111;
memory[2515]=8'b11111111;
memory[2516]=8'b11111111;
memory[2517]=8'b11111111;
memory[2518]=8'b11111111;
memory[2519]=8'b11111111;
memory[2520]=8'b11111111;
memory[2521]=8'b11111111;
memory[2522]=8'b11111111;
memory[2523]=8'b11111111;
memory[2524]=8'b11111111;
memory[2525]=8'b11111111;
memory[2526]=8'b11111111;
memory[2527]=8'b11111111;
memory[2528]=8'b11111111;
memory[2529]=8'b11111111;
memory[2530]=8'b11111111;
memory[2531]=8'b11111111;
memory[2532]=8'b11111111;
memory[2533]=8'b11111111;
memory[2534]=8'b11111111;
memory[2535]=8'b11111111;
memory[2536]=8'b11111111;
memory[2537]=8'b11111111;
memory[2538]=8'b11100000;
memory[2539]=8'b00000011;
memory[2540]=8'b11111111;
memory[2541]=8'b11111111;
memory[2542]=8'b11111111;
memory[2543]=8'b11111111;
memory[2544]=8'b11111000;
memory[2545]=8'b00000000;
memory[2546]=8'b00000000;
memory[2547]=8'b00000000;
memory[2548]=8'b00000000;
memory[2549]=8'b00000000;
memory[2550]=8'b00001111;
memory[2551]=8'b11111111;
memory[2552]=8'b11111111;
memory[2553]=8'b11111111;
memory[2554]=8'b11111111;
memory[2555]=8'b11111111;
memory[2556]=8'b11111111;
memory[2557]=8'b11111111;
memory[2558]=8'b11111111;
memory[2559]=8'b11111111;
memory[2560]=8'b11111111;
memory[2561]=8'b11111111;
memory[2562]=8'b11111111;
memory[2563]=8'b11111111;
memory[2564]=8'b11111111;
memory[2565]=8'b11111111;
memory[2566]=8'b11111111;
memory[2567]=8'b11111111;
memory[2568]=8'b11111111;
memory[2569]=8'b11111111;
memory[2570]=8'b11111111;
memory[2571]=8'b11111111;
memory[2572]=8'b11111111;
memory[2573]=8'b11111111;
memory[2574]=8'b11111111;
memory[2575]=8'b11111111;
memory[2576]=8'b11111111;
memory[2577]=8'b11111111;
memory[2578]=8'b11110000;
memory[2579]=8'b00000001;
memory[2580]=8'b11111111;
memory[2581]=8'b11111111;
memory[2582]=8'b11111111;
memory[2583]=8'b11111111;
memory[2584]=8'b11000000;
memory[2585]=8'b00000000;
memory[2586]=8'b00000000;
memory[2587]=8'b00000000;
memory[2588]=8'b00000000;
memory[2589]=8'b00000000;
memory[2590]=8'b00000000;
memory[2591]=8'b11111111;
memory[2592]=8'b11111111;
memory[2593]=8'b11111111;
memory[2594]=8'b11111111;
memory[2595]=8'b11111111;
memory[2596]=8'b11111111;
memory[2597]=8'b11111111;
memory[2598]=8'b11111111;
memory[2599]=8'b11111111;
memory[2600]=8'b11111111;
memory[2601]=8'b11111111;
memory[2602]=8'b11111111;
memory[2603]=8'b11111111;
memory[2604]=8'b11111111;
memory[2605]=8'b11111111;
memory[2606]=8'b11111111;
memory[2607]=8'b11111111;
memory[2608]=8'b11111111;
memory[2609]=8'b11111111;
memory[2610]=8'b11111111;
memory[2611]=8'b11111111;
memory[2612]=8'b11111111;
memory[2613]=8'b11111111;
memory[2614]=8'b11111111;
memory[2615]=8'b11111111;
memory[2616]=8'b11111111;
memory[2617]=8'b11111111;
memory[2618]=8'b11111000;
memory[2619]=8'b00000000;
memory[2620]=8'b11111111;
memory[2621]=8'b11111111;
memory[2622]=8'b11111111;
memory[2623]=8'b11111111;
memory[2624]=8'b11000111;
memory[2625]=8'b11000000;
memory[2626]=8'b00000000;
memory[2627]=8'b00000000;
memory[2628]=8'b00011100;
memory[2629]=8'b00000000;
memory[2630]=8'b00000000;
memory[2631]=8'b00111111;
memory[2632]=8'b11111111;
memory[2633]=8'b11111111;
memory[2634]=8'b11111111;
memory[2635]=8'b11111111;
memory[2636]=8'b11111111;
memory[2637]=8'b11111111;
memory[2638]=8'b11111111;
memory[2639]=8'b11111111;
memory[2640]=8'b11111111;
memory[2641]=8'b11111111;
memory[2642]=8'b11111111;
memory[2643]=8'b11111111;
memory[2644]=8'b11111111;
memory[2645]=8'b11111111;
memory[2646]=8'b11111111;
memory[2647]=8'b11111111;
memory[2648]=8'b11111111;
memory[2649]=8'b11111111;
memory[2650]=8'b11111111;
memory[2651]=8'b11111111;
memory[2652]=8'b11111111;
memory[2653]=8'b11111111;
memory[2654]=8'b11111111;
memory[2655]=8'b11111111;
memory[2656]=8'b11111111;
memory[2657]=8'b11111111;
memory[2658]=8'b11111100;
memory[2659]=8'b00000000;
memory[2660]=8'b01111111;
memory[2661]=8'b11111111;
memory[2662]=8'b11111111;
memory[2663]=8'b11111111;
memory[2664]=8'b11111111;
memory[2665]=8'b11111110;
memory[2666]=8'b00000000;
memory[2667]=8'b01111111;
memory[2668]=8'b11111111;
memory[2669]=8'b11111111;
memory[2670]=8'b11111111;
memory[2671]=8'b11111111;
memory[2672]=8'b11111111;
memory[2673]=8'b11111111;
memory[2674]=8'b11111111;
memory[2675]=8'b11111111;
memory[2676]=8'b11111111;
memory[2677]=8'b11111111;
memory[2678]=8'b11111111;
memory[2679]=8'b11111111;
memory[2680]=8'b11111111;
memory[2681]=8'b11111111;
memory[2682]=8'b11111111;
memory[2683]=8'b11111111;
memory[2684]=8'b11111111;
memory[2685]=8'b11111111;
memory[2686]=8'b11111111;
memory[2687]=8'b11111111;
memory[2688]=8'b11111111;
memory[2689]=8'b11111111;
memory[2690]=8'b11111111;
memory[2691]=8'b11111111;
memory[2692]=8'b11111111;
memory[2693]=8'b11111111;
memory[2694]=8'b11111111;
memory[2695]=8'b11111111;
memory[2696]=8'b11111111;
memory[2697]=8'b11111111;
memory[2698]=8'b11111110;
memory[2699]=8'b00000000;
memory[2700]=8'b00111111;
memory[2701]=8'b11111111;
memory[2702]=8'b11111111;
memory[2703]=8'b11111111;
memory[2704]=8'b11111111;
memory[2705]=8'b11111111;
memory[2706]=8'b11111111;
memory[2707]=8'b11111111;
memory[2708]=8'b11111111;
memory[2709]=8'b11111111;
memory[2710]=8'b11111111;
memory[2711]=8'b11111111;
memory[2712]=8'b11111111;
memory[2713]=8'b11111111;
memory[2714]=8'b11111111;
memory[2715]=8'b11111111;
memory[2716]=8'b11111111;
memory[2717]=8'b11111111;
memory[2718]=8'b11111111;
memory[2719]=8'b11111111;
memory[2720]=8'b11111111;
memory[2721]=8'b11111111;
memory[2722]=8'b11111111;
memory[2723]=8'b11111111;
memory[2724]=8'b11111111;
memory[2725]=8'b11111111;
memory[2726]=8'b11111111;
memory[2727]=8'b11111111;
memory[2728]=8'b11111111;
memory[2729]=8'b11111111;
memory[2730]=8'b11111111;
memory[2731]=8'b11111111;
memory[2732]=8'b11111111;
memory[2733]=8'b11111111;
memory[2734]=8'b11111111;
memory[2735]=8'b11111111;
memory[2736]=8'b11111111;
memory[2737]=8'b11111111;
memory[2738]=8'b11111111;
memory[2739]=8'b00000000;
memory[2740]=8'b00011111;
memory[2741]=8'b11111111;
memory[2742]=8'b11111111;
memory[2743]=8'b11111111;
memory[2744]=8'b11111111;
memory[2745]=8'b11111111;
memory[2746]=8'b11111111;
memory[2747]=8'b11111111;
memory[2748]=8'b11111111;
memory[2749]=8'b11111111;
memory[2750]=8'b11111111;
memory[2751]=8'b11111111;
memory[2752]=8'b11111111;
memory[2753]=8'b11111111;
memory[2754]=8'b11111111;
memory[2755]=8'b11111111;
memory[2756]=8'b11111111;
memory[2757]=8'b11111111;
memory[2758]=8'b11111111;
memory[2759]=8'b11111111;
memory[2760]=8'b11111111;
memory[2761]=8'b11111111;
memory[2762]=8'b11111111;
memory[2763]=8'b11111111;
memory[2764]=8'b11111111;
memory[2765]=8'b11111111;
memory[2766]=8'b11111111;
memory[2767]=8'b11111111;
memory[2768]=8'b11111111;
memory[2769]=8'b11111111;
memory[2770]=8'b11111111;
memory[2771]=8'b11111111;
memory[2772]=8'b11111111;
memory[2773]=8'b11111111;
memory[2774]=8'b11000000;
memory[2775]=8'b00011111;
memory[2776]=8'b11111111;
memory[2777]=8'b11111111;
memory[2778]=8'b11111111;
memory[2779]=8'b11000000;
memory[2780]=8'b00011111;
memory[2781]=8'b11111111;
memory[2782]=8'b11111111;
memory[2783]=8'b11111111;
memory[2784]=8'b11111111;
memory[2785]=8'b11111111;
memory[2786]=8'b11111111;
memory[2787]=8'b11111111;
memory[2788]=8'b11110000;
memory[2789]=8'b00000000;
memory[2790]=8'b00000000;
memory[2791]=8'b00000000;
memory[2792]=8'b00111111;
memory[2793]=8'b11111111;
memory[2794]=8'b11111111;
memory[2795]=8'b11111111;
memory[2796]=8'b11111111;
memory[2797]=8'b11111111;
memory[2798]=8'b11111111;
memory[2799]=8'b11111111;
memory[2800]=8'b11111111;
memory[2801]=8'b11111111;
memory[2802]=8'b11111111;
memory[2803]=8'b11111111;
memory[2804]=8'b11111111;
memory[2805]=8'b11111111;
memory[2806]=8'b11111111;
memory[2807]=8'b11111111;
memory[2808]=8'b11111111;
memory[2809]=8'b11111111;
memory[2810]=8'b11111111;
memory[2811]=8'b11111111;
memory[2812]=8'b11111111;
memory[2813]=8'b10000000;
memory[2814]=8'b00000000;
memory[2815]=8'b00000000;
memory[2816]=8'b00111111;
memory[2817]=8'b11111111;
memory[2818]=8'b11111111;
memory[2819]=8'b11000000;
memory[2820]=8'b00001111;
memory[2821]=8'b11111111;
memory[2822]=8'b11111111;
memory[2823]=8'b11111111;
memory[2824]=8'b11111111;
memory[2825]=8'b11111111;
memory[2826]=8'b11111111;
memory[2827]=8'b11111111;
memory[2828]=8'b11111111;
memory[2829]=8'b11100000;
memory[2830]=8'b00000011;
memory[2831]=8'b11111111;
memory[2832]=8'b11111111;
memory[2833]=8'b11111111;
memory[2834]=8'b11111111;
memory[2835]=8'b11111111;
memory[2836]=8'b11111111;
memory[2837]=8'b11111111;
memory[2838]=8'b11111111;
memory[2839]=8'b11111111;
memory[2840]=8'b11111111;
memory[2841]=8'b11111111;
memory[2842]=8'b11111111;
memory[2843]=8'b11111111;
memory[2844]=8'b11111111;
memory[2845]=8'b11111111;
memory[2846]=8'b11111111;
memory[2847]=8'b11111111;
memory[2848]=8'b11111111;
memory[2849]=8'b11111111;
memory[2850]=8'b11111111;
memory[2851]=8'b11111111;
memory[2852]=8'b11111111;
memory[2853]=8'b11111111;
memory[2854]=8'b11111000;
memory[2855]=8'b00000000;
memory[2856]=8'b00000111;
memory[2857]=8'b11111111;
memory[2858]=8'b11111111;
memory[2859]=8'b11100000;
memory[2860]=8'b00000111;
memory[2861]=8'b11111111;
memory[2862]=8'b11111111;
memory[2863]=8'b11111111;
memory[2864]=8'b11111111;
memory[2865]=8'b11111111;
memory[2866]=8'b11110111;
memory[2867]=8'b11111110;
memory[2868]=8'b00001100;
memory[2869]=8'b00000000;
memory[2870]=8'b00000001;
memory[2871]=8'b11111111;
memory[2872]=8'b11111111;
memory[2873]=8'b11111111;
memory[2874]=8'b11111111;
memory[2875]=8'b11111111;
memory[2876]=8'b11111111;
memory[2877]=8'b11111111;
memory[2878]=8'b11111111;
memory[2879]=8'b11111111;
memory[2880]=8'b11111111;
memory[2881]=8'b11111111;
memory[2882]=8'b11111111;
memory[2883]=8'b11111111;
memory[2884]=8'b11111111;
memory[2885]=8'b11111111;
memory[2886]=8'b11111111;
memory[2887]=8'b11111111;
memory[2888]=8'b11111111;
memory[2889]=8'b11111111;
memory[2890]=8'b11111111;
memory[2891]=8'b11111100;
memory[2892]=8'b00011111;
memory[2893]=8'b11111111;
memory[2894]=8'b11111111;
memory[2895]=8'b11000000;
memory[2896]=8'b00000000;
memory[2897]=8'b11111111;
memory[2898]=8'b11111111;
memory[2899]=8'b11110000;
memory[2900]=8'b00000011;
memory[2901]=8'b11111111;
memory[2902]=8'b11111111;
memory[2903]=8'b11111111;
memory[2904]=8'b11111111;
memory[2905]=8'b11111111;
memory[2906]=8'b11111111;
memory[2907]=8'b11111111;
memory[2908]=8'b11110000;
memory[2909]=8'b00000000;
memory[2910]=8'b00000001;
memory[2911]=8'b11111111;
memory[2912]=8'b11111111;
memory[2913]=8'b11111111;
memory[2914]=8'b11111111;
memory[2915]=8'b11111111;
memory[2916]=8'b11111111;
memory[2917]=8'b11111111;
memory[2918]=8'b11111111;
memory[2919]=8'b11111111;
memory[2920]=8'b11111111;
memory[2921]=8'b11111111;
memory[2922]=8'b11111111;
memory[2923]=8'b11111111;
memory[2924]=8'b11111111;
memory[2925]=8'b11111111;
memory[2926]=8'b11111111;
memory[2927]=8'b11111111;
memory[2928]=8'b11111111;
memory[2929]=8'b11111111;
memory[2930]=8'b11111111;
memory[2931]=8'b11100000;
memory[2932]=8'b11111111;
memory[2933]=8'b11111111;
memory[2934]=8'b11111110;
memory[2935]=8'b00000000;
memory[2936]=8'b00000000;
memory[2937]=8'b00111111;
memory[2938]=8'b11111111;
memory[2939]=8'b11111000;
memory[2940]=8'b00000011;
memory[2941]=8'b11111111;
memory[2942]=8'b11111111;
memory[2943]=8'b11111111;
memory[2944]=8'b11111111;
memory[2945]=8'b11111111;
memory[2946]=8'b11111111;
memory[2947]=8'b11111111;
memory[2948]=8'b11110000;
memory[2949]=8'b00000000;
memory[2950]=8'b00000111;
memory[2951]=8'b11111111;
memory[2952]=8'b11111111;
memory[2953]=8'b11111111;
memory[2954]=8'b11111111;
memory[2955]=8'b11111111;
memory[2956]=8'b11111111;
memory[2957]=8'b11111111;
memory[2958]=8'b11111111;
memory[2959]=8'b11111111;
memory[2960]=8'b11111111;
memory[2961]=8'b11111111;
memory[2962]=8'b11111111;
memory[2963]=8'b11111111;
memory[2964]=8'b11111111;
memory[2965]=8'b11111111;
memory[2966]=8'b11111111;
memory[2967]=8'b11111111;
memory[2968]=8'b11111111;
memory[2969]=8'b11111111;
memory[2970]=8'b11111111;
memory[2971]=8'b00000111;
memory[2972]=8'b11111111;
memory[2973]=8'b11111111;
memory[2974]=8'b11111111;
memory[2975]=8'b11110000;
memory[2976]=8'b00000000;
memory[2977]=8'b00001111;
memory[2978]=8'b11111111;
memory[2979]=8'b11111100;
memory[2980]=8'b00000001;
memory[2981]=8'b11111111;
memory[2982]=8'b11111111;
memory[2983]=8'b11110000;
memory[2984]=8'b11111111;
memory[2985]=8'b11111111;
memory[2986]=8'b11110000;
memory[2987]=8'b00000000;
memory[2988]=8'b00000000;
memory[2989]=8'b00000000;
memory[2990]=8'b00000000;
memory[2991]=8'b00000000;
memory[2992]=8'b00001111;
memory[2993]=8'b11111111;
memory[2994]=8'b11111111;
memory[2995]=8'b11111111;
memory[2996]=8'b11111111;
memory[2997]=8'b11111111;
memory[2998]=8'b11111111;
memory[2999]=8'b11111111;
memory[3000]=8'b11111111;
memory[3001]=8'b11111111;
memory[3002]=8'b11111111;
memory[3003]=8'b11111111;
memory[3004]=8'b11111111;
memory[3005]=8'b11111111;
memory[3006]=8'b11111111;
memory[3007]=8'b11111111;
memory[3008]=8'b11111111;
memory[3009]=8'b11111111;
memory[3010]=8'b11111000;
memory[3011]=8'b00011111;
memory[3012]=8'b11111111;
memory[3013]=8'b11110111;
memory[3014]=8'b11111111;
memory[3015]=8'b11111100;
memory[3016]=8'b00000000;
memory[3017]=8'b00000111;
memory[3018]=8'b11111111;
memory[3019]=8'b11111100;
memory[3020]=8'b00000000;
memory[3021]=8'b11111111;
memory[3022]=8'b11111110;
memory[3023]=8'b00000000;
memory[3024]=8'b00001111;
memory[3025]=8'b11111111;
memory[3026]=8'b11111111;
memory[3027]=8'b11111111;
memory[3028]=8'b00000000;
memory[3029]=8'b00000000;
memory[3030]=8'b00000111;
memory[3031]=8'b11111111;
memory[3032]=8'b11111111;
memory[3033]=8'b11111111;
memory[3034]=8'b11111111;
memory[3035]=8'b11111111;
memory[3036]=8'b11111111;
memory[3037]=8'b11111111;
memory[3038]=8'b11111111;
memory[3039]=8'b11111111;
memory[3040]=8'b11111111;
memory[3041]=8'b11111111;
memory[3042]=8'b11111111;
memory[3043]=8'b11111111;
memory[3044]=8'b11111111;
memory[3045]=8'b11111111;
memory[3046]=8'b11111111;
memory[3047]=8'b11111111;
memory[3048]=8'b11111111;
memory[3049]=8'b11111111;
memory[3050]=8'b11110001;
memory[3051]=8'b11111111;
memory[3052]=8'b11111111;
memory[3053]=8'b11001111;
memory[3054]=8'b11111111;
memory[3055]=8'b11111110;
memory[3056]=8'b00000000;
memory[3057]=8'b00000011;
memory[3058]=8'b11111111;
memory[3059]=8'b11111110;
memory[3060]=8'b00000000;
memory[3061]=8'b11111111;
memory[3062]=8'b11111100;
memory[3063]=8'b00000000;
memory[3064]=8'b00000011;
memory[3065]=8'b11111111;
memory[3066]=8'b11111111;
memory[3067]=8'b11111111;
memory[3068]=8'b11110000;
memory[3069]=8'b00000000;
memory[3070]=8'b00000011;
memory[3071]=8'b11111111;
memory[3072]=8'b11111111;
memory[3073]=8'b11111111;
memory[3074]=8'b11111111;
memory[3075]=8'b11111111;
memory[3076]=8'b11111111;
memory[3077]=8'b11111111;
memory[3078]=8'b11111111;
memory[3079]=8'b11111111;
memory[3080]=8'b11111111;
memory[3081]=8'b11111111;
memory[3082]=8'b11111111;
memory[3083]=8'b11111111;
memory[3084]=8'b11111111;
memory[3085]=8'b11111111;
memory[3086]=8'b11111111;
memory[3087]=8'b11111111;
memory[3088]=8'b11111111;
memory[3089]=8'b11111111;
memory[3090]=8'b11001111;
memory[3091]=8'b11111111;
memory[3092]=8'b11111111;
memory[3093]=8'b10001111;
memory[3094]=8'b11011111;
memory[3095]=8'b11111110;
memory[3096]=8'b00000000;
memory[3097]=8'b00000001;
memory[3098]=8'b11111111;
memory[3099]=8'b11111111;
memory[3100]=8'b00000000;
memory[3101]=8'b01111111;
memory[3102]=8'b11111100;
memory[3103]=8'b00111100;
memory[3104]=8'b00000001;
memory[3105]=8'b11111111;
memory[3106]=8'b11110000;
memory[3107]=8'b00001111;
memory[3108]=8'b11100000;
memory[3109]=8'b00000000;
memory[3110]=8'b01111111;
memory[3111]=8'b11111111;
memory[3112]=8'b11111111;
memory[3113]=8'b11111111;
memory[3114]=8'b11111111;
memory[3115]=8'b11111111;
memory[3116]=8'b11111111;
memory[3117]=8'b11111111;
memory[3118]=8'b11111111;
memory[3119]=8'b11111111;
memory[3120]=8'b11111111;
memory[3121]=8'b11111111;
memory[3122]=8'b11111111;
memory[3123]=8'b11111111;
memory[3124]=8'b11111111;
memory[3125]=8'b11111111;
memory[3126]=8'b11111111;
memory[3127]=8'b11111111;
memory[3128]=8'b11111111;
memory[3129]=8'b11111111;
memory[3130]=8'b00111111;
memory[3131]=8'b11111111;
memory[3132]=8'b11111111;
memory[3133]=8'b10001111;
memory[3134]=8'b00011111;
memory[3135]=8'b11111100;
memory[3136]=8'b00000000;
memory[3137]=8'b00000000;
memory[3138]=8'b11111111;
memory[3139]=8'b11111111;
memory[3140]=8'b00000000;
memory[3141]=8'b01111111;
memory[3142]=8'b11111111;
memory[3143]=8'b11111110;
memory[3144]=8'b00000000;
memory[3145]=8'b11111111;
memory[3146]=8'b11110000;
memory[3147]=8'b00111111;
memory[3148]=8'b11111100;
memory[3149]=8'b00000011;
memory[3150]=8'b11111111;
memory[3151]=8'b11111111;
memory[3152]=8'b11111111;
memory[3153]=8'b11111111;
memory[3154]=8'b11111111;
memory[3155]=8'b11111111;
memory[3156]=8'b11111111;
memory[3157]=8'b11111111;
memory[3158]=8'b11111111;
memory[3159]=8'b11111111;
memory[3160]=8'b11111111;
memory[3161]=8'b11111111;
memory[3162]=8'b11111111;
memory[3163]=8'b11111111;
memory[3164]=8'b11111111;
memory[3165]=8'b11111111;
memory[3166]=8'b11111111;
memory[3167]=8'b11111111;
memory[3168]=8'b11111111;
memory[3169]=8'b11111111;
memory[3170]=8'b11111111;
memory[3171]=8'b11110111;
memory[3172]=8'b11111111;
memory[3173]=8'b10000000;
memory[3174]=8'b00111111;
memory[3175]=8'b11110000;
memory[3176]=8'b00000000;
memory[3177]=8'b00000000;
memory[3178]=8'b01111111;
memory[3179]=8'b11111111;
memory[3180]=8'b00000000;
memory[3181]=8'b01111111;
memory[3182]=8'b11111111;
memory[3183]=8'b11111000;
memory[3184]=8'b00000000;
memory[3185]=8'b01111111;
memory[3186]=8'b11111111;
memory[3187]=8'b11111111;
memory[3188]=8'b11111110;
memory[3189]=8'b00000001;
memory[3190]=8'b11111111;
memory[3191]=8'b11111111;
memory[3192]=8'b11111111;
memory[3193]=8'b11111111;
memory[3194]=8'b11111111;
memory[3195]=8'b11111111;
memory[3196]=8'b11111111;
memory[3197]=8'b11111111;
memory[3198]=8'b11111111;
memory[3199]=8'b11111111;
memory[3200]=8'b11111111;
memory[3201]=8'b11111111;
memory[3202]=8'b11111111;
memory[3203]=8'b11111111;
memory[3204]=8'b11111111;
memory[3205]=8'b11111111;
memory[3206]=8'b11111111;
memory[3207]=8'b11111111;
memory[3208]=8'b11111111;
memory[3209]=8'b11111111;
memory[3210]=8'b11111111;
memory[3211]=8'b11101111;
memory[3212]=8'b11111111;
memory[3213]=8'b10000000;
memory[3214]=8'b00111111;
memory[3215]=8'b11111111;
memory[3216]=8'b00000000;
memory[3217]=8'b00000000;
memory[3218]=8'b00111111;
memory[3219]=8'b11111111;
memory[3220]=8'b00000000;
memory[3221]=8'b00111111;
memory[3222]=8'b11111111;
memory[3223]=8'b11100000;
memory[3224]=8'b00000000;
memory[3225]=8'b00111111;
memory[3226]=8'b11111111;
memory[3227]=8'b11110000;
memory[3228]=8'b00000000;
memory[3229]=8'b00000000;
memory[3230]=8'b00000000;
memory[3231]=8'b00111111;
memory[3232]=8'b11111111;
memory[3233]=8'b11111111;
memory[3234]=8'b11111111;
memory[3235]=8'b11111111;
memory[3236]=8'b11111111;
memory[3237]=8'b11111111;
memory[3238]=8'b11111111;
memory[3239]=8'b11111111;
memory[3240]=8'b11111111;
memory[3241]=8'b11111111;
memory[3242]=8'b11111111;
memory[3243]=8'b11111111;
memory[3244]=8'b11111111;
memory[3245]=8'b11111111;
memory[3246]=8'b11111111;
memory[3247]=8'b11111111;
memory[3248]=8'b11111111;
memory[3249]=8'b11111111;
memory[3250]=8'b11111111;
memory[3251]=8'b11001111;
memory[3252]=8'b11111001;
memory[3253]=8'b00000000;
memory[3254]=8'b00001111;
memory[3255]=8'b11111111;
memory[3256]=8'b10000000;
memory[3257]=8'b00000000;
memory[3258]=8'b00111111;
memory[3259]=8'b11111111;
memory[3260]=8'b10000000;
memory[3261]=8'b00111111;
memory[3262]=8'b11111111;
memory[3263]=8'b10000000;
memory[3264]=8'b00000000;
memory[3265]=8'b00111111;
memory[3266]=8'b11111111;
memory[3267]=8'b11111000;
memory[3268]=8'b00000001;
memory[3269]=8'b11111111;
memory[3270]=8'b11111111;
memory[3271]=8'b11111111;
memory[3272]=8'b11111111;
memory[3273]=8'b11111111;
memory[3274]=8'b11111111;
memory[3275]=8'b11111111;
memory[3276]=8'b11111111;
memory[3277]=8'b11111111;
memory[3278]=8'b11111111;
memory[3279]=8'b11111111;
memory[3280]=8'b11111111;
memory[3281]=8'b11111111;
memory[3282]=8'b11111111;
memory[3283]=8'b11111111;
memory[3284]=8'b11111111;
memory[3285]=8'b11111111;
memory[3286]=8'b11111111;
memory[3287]=8'b11111111;
memory[3288]=8'b11111111;
memory[3289]=8'b11101111;
memory[3290]=8'b11100111;
memory[3291]=8'b10011111;
memory[3292]=8'b11100000;
memory[3293]=8'b00000000;
memory[3294]=8'b00001111;
memory[3295]=8'b11111100;
memory[3296]=8'b00000000;
memory[3297]=8'b00000000;
memory[3298]=8'b00011111;
memory[3299]=8'b11111111;
memory[3300]=8'b10000000;
memory[3301]=8'b00111111;
memory[3302]=8'b11111111;
memory[3303]=8'b11111111;
memory[3304]=8'b11000000;
memory[3305]=8'b00011111;
memory[3306]=8'b11111111;
memory[3307]=8'b11111111;
memory[3308]=8'b11101111;
memory[3309]=8'b11111111;
memory[3310]=8'b11111111;
memory[3311]=8'b11111111;
memory[3312]=8'b11111111;
memory[3313]=8'b11111111;
memory[3314]=8'b11111111;
memory[3315]=8'b11111111;
memory[3316]=8'b11111111;
memory[3317]=8'b11111111;
memory[3318]=8'b11111111;
memory[3319]=8'b11111111;
memory[3320]=8'b11111111;
memory[3321]=8'b11111111;
memory[3322]=8'b11111111;
memory[3323]=8'b11111111;
memory[3324]=8'b11111111;
memory[3325]=8'b11111111;
memory[3326]=8'b11111111;
memory[3327]=8'b11111111;
memory[3328]=8'b11111111;
memory[3329]=8'b10001111;
memory[3330]=8'b11001111;
memory[3331]=8'b00011111;
memory[3332]=8'b00000000;
memory[3333]=8'b00000000;
memory[3334]=8'b00000011;
memory[3335]=8'b11110000;
memory[3336]=8'b00000000;
memory[3337]=8'b00000000;
memory[3338]=8'b00001111;
memory[3339]=8'b11111111;
memory[3340]=8'b00000000;
memory[3341]=8'b00111110;
memory[3342]=8'b01111111;
memory[3343]=8'b11111111;
memory[3344]=8'b11100000;
memory[3345]=8'b00011111;
memory[3346]=8'b11111111;
memory[3347]=8'b11111111;
memory[3348]=8'b11111111;
memory[3349]=8'b11111111;
memory[3350]=8'b11111111;
memory[3351]=8'b11111111;
memory[3352]=8'b11111111;
memory[3353]=8'b11111111;
memory[3354]=8'b11111111;
memory[3355]=8'b11111111;
memory[3356]=8'b11111111;
memory[3357]=8'b11111111;
memory[3358]=8'b11111111;
memory[3359]=8'b11111111;
memory[3360]=8'b11111111;
memory[3361]=8'b11111111;
memory[3362]=8'b11111111;
memory[3363]=8'b11111111;
memory[3364]=8'b11111111;
memory[3365]=8'b11111111;
memory[3366]=8'b11111111;
memory[3367]=8'b11111111;
memory[3368]=8'b11111111;
memory[3369]=8'b00011111;
memory[3370]=8'b11000110;
memory[3371]=8'b00111110;
memory[3372]=8'b00000000;
memory[3373]=8'b00000000;
memory[3374]=8'b00000111;
memory[3375]=8'b11110000;
memory[3376]=8'b00000000;
memory[3377]=8'b00000000;
memory[3378]=8'b00001111;
memory[3379]=8'b11111111;
memory[3380]=8'b00000000;
memory[3381]=8'b00111100;
memory[3382]=8'b00011111;
memory[3383]=8'b11111111;
memory[3384]=8'b11100000;
memory[3385]=8'b00011111;
memory[3386]=8'b11111111;
memory[3387]=8'b11111111;
memory[3388]=8'b11111111;
memory[3389]=8'b11111111;
memory[3390]=8'b11111111;
memory[3391]=8'b11111111;
memory[3392]=8'b11111111;
memory[3393]=8'b11111111;
memory[3394]=8'b11111111;
memory[3395]=8'b11111111;
memory[3396]=8'b11111111;
memory[3397]=8'b11111111;
memory[3398]=8'b11111111;
memory[3399]=8'b11111111;
memory[3400]=8'b11111111;
memory[3401]=8'b11111111;
memory[3402]=8'b11111111;
memory[3403]=8'b11111111;
memory[3404]=8'b11111111;
memory[3405]=8'b11111111;
memory[3406]=8'b11111111;
memory[3407]=8'b11111111;
memory[3408]=8'b11111110;
memory[3409]=8'b00001111;
memory[3410]=8'b11000000;
memory[3411]=8'b00111100;
memory[3412]=8'b00000000;
memory[3413]=8'b00000000;
memory[3414]=8'b00001111;
memory[3415]=8'b11110000;
memory[3416]=8'b00000000;
memory[3417]=8'b00000000;
memory[3418]=8'b00000111;
memory[3419]=8'b11111111;
memory[3420]=8'b00000000;
memory[3421]=8'b00111100;
memory[3422]=8'b00011111;
memory[3423]=8'b11111111;
memory[3424]=8'b11100000;
memory[3425]=8'b00011111;
memory[3426]=8'b11111111;
memory[3427]=8'b11111111;
memory[3428]=8'b11111111;
memory[3429]=8'b11111111;
memory[3430]=8'b11111111;
memory[3431]=8'b11111111;
memory[3432]=8'b11111111;
memory[3433]=8'b11111111;
memory[3434]=8'b11111111;
memory[3435]=8'b11111111;
memory[3436]=8'b11111111;
memory[3437]=8'b11111111;
memory[3438]=8'b11111111;
memory[3439]=8'b11111111;
memory[3440]=8'b11111111;
memory[3441]=8'b11111111;
memory[3442]=8'b11111111;
memory[3443]=8'b11111111;
memory[3444]=8'b11111111;
memory[3445]=8'b11111111;
memory[3446]=8'b11111111;
memory[3447]=8'b11111111;
memory[3448]=8'b11111000;
memory[3449]=8'b00000011;
memory[3450]=8'b11000000;
memory[3451]=8'b00011000;
memory[3452]=8'b00000000;
memory[3453]=8'b00000000;
memory[3454]=8'b11111111;
memory[3455]=8'b11110000;
memory[3456]=8'b00000000;
memory[3457]=8'b00000000;
memory[3458]=8'b00000111;
memory[3459]=8'b11111110;
memory[3460]=8'b00000000;
memory[3461]=8'b00111110;
memory[3462]=8'b00111111;
memory[3463]=8'b11111111;
memory[3464]=8'b11100000;
memory[3465]=8'b00111111;
memory[3466]=8'b11111111;
memory[3467]=8'b11111111;
memory[3468]=8'b11111111;
memory[3469]=8'b11111111;
memory[3470]=8'b11111111;
memory[3471]=8'b11111111;
memory[3472]=8'b11111111;
memory[3473]=8'b11111111;
memory[3474]=8'b11111111;
memory[3475]=8'b11111111;
memory[3476]=8'b11111111;
memory[3477]=8'b11111111;
memory[3478]=8'b11111111;
memory[3479]=8'b11111111;
memory[3480]=8'b11111111;
memory[3481]=8'b11111111;
memory[3482]=8'b11111111;
memory[3483]=8'b11111111;
memory[3484]=8'b11111111;
memory[3485]=8'b11111111;
memory[3486]=8'b11111111;
memory[3487]=8'b11111111;
memory[3488]=8'b11110000;
memory[3489]=8'b00000011;
memory[3490]=8'b00000000;
memory[3491]=8'b00000000;
memory[3492]=8'b00000000;
memory[3493]=8'b00000111;
memory[3494]=8'b11111111;
memory[3495]=8'b11110000;
memory[3496]=8'b00000000;
memory[3497]=8'b00000000;
memory[3498]=8'b00000111;
memory[3499]=8'b11111110;
memory[3500]=8'b00000000;
memory[3501]=8'b00011110;
memory[3502]=8'b00111111;
memory[3503]=8'b11111111;
memory[3504]=8'b11000000;
memory[3505]=8'b00111111;
memory[3506]=8'b11111111;
memory[3507]=8'b11111111;
memory[3508]=8'b11111111;
memory[3509]=8'b11111111;
memory[3510]=8'b11111111;
memory[3511]=8'b11111111;
memory[3512]=8'b11111111;
memory[3513]=8'b11111111;
memory[3514]=8'b11111111;
memory[3515]=8'b11111111;
memory[3516]=8'b11111111;
memory[3517]=8'b11111111;
memory[3518]=8'b11111111;
memory[3519]=8'b11111111;
memory[3520]=8'b11111111;
memory[3521]=8'b11111111;
memory[3522]=8'b11111111;
memory[3523]=8'b11111111;
memory[3524]=8'b11111111;
memory[3525]=8'b11111111;
memory[3526]=8'b11111111;
memory[3527]=8'b11111111;
memory[3528]=8'b11000000;
memory[3529]=8'b00000000;
memory[3530]=8'b00000000;
memory[3531]=8'b00000000;
memory[3532]=8'b00000000;
memory[3533]=8'b11111111;
memory[3534]=8'b11110000;
memory[3535]=8'b00000000;
memory[3536]=8'b00000000;
memory[3537]=8'b00000000;
memory[3538]=8'b00000001;
memory[3539]=8'b11111000;
memory[3540]=8'b00000000;
memory[3541]=8'b00011110;
memory[3542]=8'b01111111;
memory[3543]=8'b11111111;
memory[3544]=8'b10000000;
memory[3545]=8'b00111111;
memory[3546]=8'b11111111;
memory[3547]=8'b11111111;
memory[3548]=8'b11111111;
memory[3549]=8'b11111111;
memory[3550]=8'b11111111;
memory[3551]=8'b11111111;
memory[3552]=8'b11111111;
memory[3553]=8'b11111111;
memory[3554]=8'b11111111;
memory[3555]=8'b11111111;
memory[3556]=8'b11111111;
memory[3557]=8'b11111111;
memory[3558]=8'b11111111;
memory[3559]=8'b11111111;
memory[3560]=8'b11111111;
memory[3561]=8'b11111111;
memory[3562]=8'b11111111;
memory[3563]=8'b11111111;
memory[3564]=8'b11111111;
memory[3565]=8'b11111111;
memory[3566]=8'b11111111;
memory[3567]=8'b11111111;
memory[3568]=8'b00000000;
memory[3569]=8'b00000000;
memory[3570]=8'b00000000;
memory[3571]=8'b00000000;
memory[3572]=8'b00111111;
memory[3573]=8'b11111111;
memory[3574]=8'b11110000;
memory[3575]=8'b00000000;
memory[3576]=8'b00000000;
memory[3577]=8'b00000000;
memory[3578]=8'b00000000;
memory[3579]=8'b00000000;
memory[3580]=8'b00000000;
memory[3581]=8'b00111111;
memory[3582]=8'b11111111;
memory[3583]=8'b11111111;
memory[3584]=8'b00000000;
memory[3585]=8'b01111111;
memory[3586]=8'b11111111;
memory[3587]=8'b11111111;
memory[3588]=8'b11111111;
memory[3589]=8'b11111111;
memory[3590]=8'b11111111;
memory[3591]=8'b11111111;
memory[3592]=8'b11111111;
memory[3593]=8'b11111111;
memory[3594]=8'b11111111;
memory[3595]=8'b11111111;
memory[3596]=8'b11111111;
memory[3597]=8'b11111111;
memory[3598]=8'b11111111;
memory[3599]=8'b11111111;
memory[3600]=8'b11111111;
memory[3601]=8'b11111111;
memory[3602]=8'b11111111;
memory[3603]=8'b11111111;
memory[3604]=8'b11111111;
memory[3605]=8'b11111111;
memory[3606]=8'b11111111;
memory[3607]=8'b11111100;
memory[3608]=8'b00000000;
memory[3609]=8'b00011100;
memory[3610]=8'b00011111;
memory[3611]=8'b11111111;
memory[3612]=8'b11111111;
memory[3613]=8'b11111111;
memory[3614]=8'b11111000;
memory[3615]=8'b00000000;
memory[3616]=8'b00000000;
memory[3617]=8'b00000000;
memory[3618]=8'b00000000;
memory[3619]=8'b00000000;
memory[3620]=8'b00000000;
memory[3621]=8'b00111111;
memory[3622]=8'b11111111;
memory[3623]=8'b11111110;
memory[3624]=8'b00000000;
memory[3625]=8'b11111111;
memory[3626]=8'b11111111;
memory[3627]=8'b11111111;
memory[3628]=8'b11111111;
memory[3629]=8'b11111111;
memory[3630]=8'b11111111;
memory[3631]=8'b11111111;
memory[3632]=8'b11111111;
memory[3633]=8'b11111111;
memory[3634]=8'b11111111;
memory[3635]=8'b11111111;
memory[3636]=8'b11111111;
memory[3637]=8'b11111111;
memory[3638]=8'b11111111;
memory[3639]=8'b11111111;
memory[3640]=8'b11111111;
memory[3641]=8'b11111111;
memory[3642]=8'b11111111;
memory[3643]=8'b11111111;
memory[3644]=8'b11111111;
memory[3645]=8'b11111111;
memory[3646]=8'b11111111;
memory[3647]=8'b11111000;
memory[3648]=8'b00000000;
memory[3649]=8'b01111100;
memory[3650]=8'b11111111;
memory[3651]=8'b11111111;
memory[3652]=8'b11111111;
memory[3653]=8'b11100111;
memory[3654]=8'b11111111;
memory[3655]=8'b00000000;
memory[3656]=8'b00000000;
memory[3657]=8'b00000000;
memory[3658]=8'b00000000;
memory[3659]=8'b00000000;
memory[3660]=8'b00000000;
memory[3661]=8'b00111111;
memory[3662]=8'b11111111;
memory[3663]=8'b11111110;
memory[3664]=8'b00000001;
memory[3665]=8'b11111111;
memory[3666]=8'b11111111;
memory[3667]=8'b11111111;
memory[3668]=8'b11111111;
memory[3669]=8'b11111111;
memory[3670]=8'b11111111;
memory[3671]=8'b11111111;
memory[3672]=8'b11111111;
memory[3673]=8'b11111111;
memory[3674]=8'b11111111;
memory[3675]=8'b11111111;
memory[3676]=8'b11111111;
memory[3677]=8'b11111111;
memory[3678]=8'b11111111;
memory[3679]=8'b11111111;
memory[3680]=8'b11111111;
memory[3681]=8'b11111111;
memory[3682]=8'b11111111;
memory[3683]=8'b11111111;
memory[3684]=8'b11111111;
memory[3685]=8'b11111111;
memory[3686]=8'b11111111;
memory[3687]=8'b11100000;
memory[3688]=8'b00000000;
memory[3689]=8'b11111111;
memory[3690]=8'b11111111;
memory[3691]=8'b11111111;
memory[3692]=8'b11111111;
memory[3693]=8'b11100001;
memory[3694]=8'b11111111;
memory[3695]=8'b10000000;
memory[3696]=8'b00000000;
memory[3697]=8'b00000000;
memory[3698]=8'b00000000;
memory[3699]=8'b00000000;
memory[3700]=8'b00000000;
memory[3701]=8'b00111111;
memory[3702]=8'b11111111;
memory[3703]=8'b11111100;
memory[3704]=8'b00000011;
memory[3705]=8'b11111111;
memory[3706]=8'b11111111;
memory[3707]=8'b11111111;
memory[3708]=8'b11111111;
memory[3709]=8'b11111111;
memory[3710]=8'b11111111;
memory[3711]=8'b11111111;
memory[3712]=8'b11111111;
memory[3713]=8'b11111111;
memory[3714]=8'b11111111;
memory[3715]=8'b11111111;
memory[3716]=8'b11111111;
memory[3717]=8'b11111111;
memory[3718]=8'b11111111;
memory[3719]=8'b11111111;
memory[3720]=8'b11111111;
memory[3721]=8'b11111111;
memory[3722]=8'b11111111;
memory[3723]=8'b11111111;
memory[3724]=8'b11111111;
memory[3725]=8'b11111111;
memory[3726]=8'b11111111;
memory[3727]=8'b11100000;
memory[3728]=8'b00000001;
memory[3729]=8'b11111111;
memory[3730]=8'b11111111;
memory[3731]=8'b11111110;
memory[3732]=8'b00111111;
memory[3733]=8'b11100000;
memory[3734]=8'b00000000;
memory[3735]=8'b00000000;
memory[3736]=8'b00000000;
memory[3737]=8'b00000000;
memory[3738]=8'b00000000;
memory[3739]=8'b00000000;
memory[3740]=8'b00000000;
memory[3741]=8'b01111111;
memory[3742]=8'b11111111;
memory[3743]=8'b11111000;
memory[3744]=8'b00000111;
memory[3745]=8'b11111111;
memory[3746]=8'b11111111;
memory[3747]=8'b11111111;
memory[3748]=8'b11111111;
memory[3749]=8'b11111111;
memory[3750]=8'b11111111;
memory[3751]=8'b11111111;
memory[3752]=8'b11111111;
memory[3753]=8'b11111111;
memory[3754]=8'b11111111;
memory[3755]=8'b11111111;
memory[3756]=8'b11111111;
memory[3757]=8'b11111111;
memory[3758]=8'b11111111;
memory[3759]=8'b11111111;
memory[3760]=8'b11111111;
memory[3761]=8'b11111111;
memory[3762]=8'b11111111;
memory[3763]=8'b11111111;
memory[3764]=8'b11111111;
memory[3765]=8'b11111111;
memory[3766]=8'b11111111;
memory[3767]=8'b11110000;
memory[3768]=8'b00000011;
memory[3769]=8'b11111111;
memory[3770]=8'b11111111;
memory[3771]=8'b11111100;
memory[3772]=8'b00000011;
memory[3773]=8'b11000000;
memory[3774]=8'b00000000;
memory[3775]=8'b00000000;
memory[3776]=8'b00000000;
memory[3777]=8'b00000000;
memory[3778]=8'b00000000;
memory[3779]=8'b00000000;
memory[3780]=8'b00000000;
memory[3781]=8'b11111111;
memory[3782]=8'b11111111;
memory[3783]=8'b11110000;
memory[3784]=8'b00001111;
memory[3785]=8'b11111111;
memory[3786]=8'b11111111;
memory[3787]=8'b11111111;
memory[3788]=8'b11111111;
memory[3789]=8'b11111111;
memory[3790]=8'b11111111;
memory[3791]=8'b11111111;
memory[3792]=8'b11111111;
memory[3793]=8'b11111111;
memory[3794]=8'b11111111;
memory[3795]=8'b11111111;
memory[3796]=8'b11111111;
memory[3797]=8'b11111111;
memory[3798]=8'b11111111;
memory[3799]=8'b11111111;
memory[3800]=8'b11111111;
memory[3801]=8'b11111111;
memory[3802]=8'b11111111;
memory[3803]=8'b11111111;
memory[3804]=8'b11111111;
memory[3805]=8'b11111111;
memory[3806]=8'b11111111;
memory[3807]=8'b11100000;
memory[3808]=8'b00001111;
memory[3809]=8'b11100000;
memory[3810]=8'b00000111;
memory[3811]=8'b11111000;
memory[3812]=8'b00000000;
memory[3813]=8'b00000000;
memory[3814]=8'b00000000;
memory[3815]=8'b00000000;
memory[3816]=8'b00000000;
memory[3817]=8'b00000000;
memory[3818]=8'b00000000;
memory[3819]=8'b00000000;
memory[3820]=8'b00000001;
memory[3821]=8'b11111111;
memory[3822]=8'b11111111;
memory[3823]=8'b11100000;
memory[3824]=8'b00011111;
memory[3825]=8'b11111111;
memory[3826]=8'b11111111;
memory[3827]=8'b11111111;
memory[3828]=8'b11111111;
memory[3829]=8'b11111111;
memory[3830]=8'b11111111;
memory[3831]=8'b11111111;
memory[3832]=8'b11111111;
memory[3833]=8'b11111111;
memory[3834]=8'b11111111;
memory[3835]=8'b11111111;
memory[3836]=8'b11111111;
memory[3837]=8'b11111111;
memory[3838]=8'b11111111;
memory[3839]=8'b11111111;
memory[3840]=8'b11111111;
memory[3841]=8'b11111111;
memory[3842]=8'b11111111;
memory[3843]=8'b11111111;
memory[3844]=8'b11111111;
memory[3845]=8'b11111111;
memory[3846]=8'b11111111;
memory[3847]=8'b11000000;
memory[3848]=8'b11111111;
memory[3849]=8'b00000000;
memory[3850]=8'b00000000;
memory[3851]=8'b00000000;
memory[3852]=8'b00000000;
memory[3853]=8'b00000000;
memory[3854]=8'b00000000;
memory[3855]=8'b00000000;
memory[3856]=8'b11111100;
memory[3857]=8'b00000000;
memory[3858]=8'b00000000;
memory[3859]=8'b00000000;
memory[3860]=8'b00000011;
memory[3861]=8'b11111111;
memory[3862]=8'b11111111;
memory[3863]=8'b10000000;
memory[3864]=8'b01111111;
memory[3865]=8'b11111111;
memory[3866]=8'b11111111;
memory[3867]=8'b11111111;
memory[3868]=8'b11111111;
memory[3869]=8'b11111111;
memory[3870]=8'b11111111;
memory[3871]=8'b11111111;
memory[3872]=8'b11111111;
memory[3873]=8'b11111111;
memory[3874]=8'b11111111;
memory[3875]=8'b11111111;
memory[3876]=8'b11111111;
memory[3877]=8'b11111111;
memory[3878]=8'b11111111;
memory[3879]=8'b11111111;
memory[3880]=8'b11111111;
memory[3881]=8'b11111111;
memory[3882]=8'b11111111;
memory[3883]=8'b11111111;
memory[3884]=8'b11111111;
memory[3885]=8'b11111111;
memory[3886]=8'b11111111;
memory[3887]=8'b10000111;
memory[3888]=8'b11111000;
memory[3889]=8'b00000011;
memory[3890]=8'b11111100;
memory[3891]=8'b00000000;
memory[3892]=8'b00000000;
memory[3893]=8'b00000000;
memory[3894]=8'b00000000;
memory[3895]=8'b00011111;
memory[3896]=8'b11111111;
memory[3897]=8'b11000000;
memory[3898]=8'b00000000;
memory[3899]=8'b00000000;
memory[3900]=8'b00011111;
memory[3901]=8'b11111111;
memory[3902]=8'b11111111;
memory[3903]=8'b00000000;
memory[3904]=8'b11111111;
memory[3905]=8'b11111111;
memory[3906]=8'b11111111;
memory[3907]=8'b11111111;
memory[3908]=8'b11111111;
memory[3909]=8'b11111111;
memory[3910]=8'b11111111;
memory[3911]=8'b11111111;
memory[3912]=8'b11111111;
memory[3913]=8'b11111111;
memory[3914]=8'b11111111;
memory[3915]=8'b11111111;
memory[3916]=8'b11111111;
memory[3917]=8'b11111111;
memory[3918]=8'b11111111;
memory[3919]=8'b11111111;
memory[3920]=8'b11111111;
memory[3921]=8'b11111111;
memory[3922]=8'b11111111;
memory[3923]=8'b11111111;
memory[3924]=8'b11111111;
memory[3925]=8'b11111111;
memory[3926]=8'b11111111;
memory[3927]=8'b11111111;
memory[3928]=8'b11000000;
memory[3929]=8'b00011111;
memory[3930]=8'b11111111;
memory[3931]=8'b11110000;
memory[3932]=8'b00000000;
memory[3933]=8'b00000000;
memory[3934]=8'b00000000;
memory[3935]=8'b11111111;
memory[3936]=8'b11111111;
memory[3937]=8'b11111110;
memory[3938]=8'b00000000;
memory[3939]=8'b00000000;
memory[3940]=8'b11111111;
memory[3941]=8'b11111111;
memory[3942]=8'b11111111;
memory[3943]=8'b00000001;
memory[3944]=8'b11111111;
memory[3945]=8'b11111111;
memory[3946]=8'b11111111;
memory[3947]=8'b11111111;
memory[3948]=8'b11111111;
memory[3949]=8'b11111111;
memory[3950]=8'b11111111;
memory[3951]=8'b11111111;
memory[3952]=8'b11111111;
memory[3953]=8'b11111111;
memory[3954]=8'b11111111;
memory[3955]=8'b11111111;
memory[3956]=8'b11111111;
memory[3957]=8'b11111111;
memory[3958]=8'b11111111;
memory[3959]=8'b11111111;
memory[3960]=8'b11111111;
memory[3961]=8'b11111111;
memory[3962]=8'b11111111;
memory[3963]=8'b11111111;
memory[3964]=8'b11111111;
memory[3965]=8'b11111111;
memory[3966]=8'b11111111;
memory[3967]=8'b11111111;
memory[3968]=8'b00000000;
memory[3969]=8'b01111110;
memory[3970]=8'b01111111;
memory[3971]=8'b11111111;
memory[3972]=8'b10000000;
memory[3973]=8'b00000000;
memory[3974]=8'b00001111;
memory[3975]=8'b11111100;
memory[3976]=8'b00000000;
memory[3977]=8'b11111111;
memory[3978]=8'b11110000;
memory[3979]=8'b00011111;
memory[3980]=8'b11111111;
memory[3981]=8'b11111111;
memory[3982]=8'b11111110;
memory[3983]=8'b00000011;
memory[3984]=8'b11111111;
memory[3985]=8'b11111111;
memory[3986]=8'b11111111;
memory[3987]=8'b11111111;
memory[3988]=8'b11111111;
memory[3989]=8'b11111111;
memory[3990]=8'b11111111;
memory[3991]=8'b11111111;
memory[3992]=8'b11111111;
memory[3993]=8'b11111111;
memory[3994]=8'b11111111;
memory[3995]=8'b11111111;
memory[3996]=8'b11111111;
memory[3997]=8'b11111111;
memory[3998]=8'b11111111;
memory[3999]=8'b11111111;
memory[4000]=8'b11111111;
memory[4001]=8'b11111111;
memory[4002]=8'b11111111;
memory[4003]=8'b11111111;
memory[4004]=8'b11111111;
memory[4005]=8'b11111111;
memory[4006]=8'b11111111;
memory[4007]=8'b11111100;
memory[4008]=8'b00000000;
memory[4009]=8'b11111111;
memory[4010]=8'b00000000;
memory[4011]=8'b01111111;
memory[4012]=8'b11111110;
memory[4013]=8'b00000000;
memory[4014]=8'b11111111;
memory[4015]=8'b10000000;
memory[4016]=8'b00111000;
memory[4017]=8'b00000111;
memory[4018]=8'b11111111;
memory[4019]=8'b11111111;
memory[4020]=8'b11111111;
memory[4021]=8'b11111111;
memory[4022]=8'b11111100;
memory[4023]=8'b00000111;
memory[4024]=8'b11111111;
memory[4025]=8'b11111111;
memory[4026]=8'b10000000;
memory[4027]=8'b00000000;
memory[4028]=8'b00111111;
memory[4029]=8'b11111111;
memory[4030]=8'b11111111;
memory[4031]=8'b11111111;
memory[4032]=8'b11111111;
memory[4033]=8'b11111111;
memory[4034]=8'b11111111;
memory[4035]=8'b11111111;
memory[4036]=8'b11111111;
memory[4037]=8'b11111111;
memory[4038]=8'b11111111;
memory[4039]=8'b11111111;
memory[4040]=8'b11111111;
memory[4041]=8'b11111111;
memory[4042]=8'b11111111;
memory[4043]=8'b11111111;
memory[4044]=8'b11111111;
memory[4045]=8'b11111111;
memory[4046]=8'b11111111;
memory[4047]=8'b11111000;
memory[4048]=8'b00000001;
memory[4049]=8'b11111111;
memory[4050]=8'b11111111;
memory[4051]=8'b11000011;
memory[4052]=8'b11111111;
memory[4053]=8'b11111111;
memory[4054]=8'b11111100;
memory[4055]=8'b00001111;
memory[4056]=8'b11111111;
memory[4057]=8'b11111111;
memory[4058]=8'b11111111;
memory[4059]=8'b11111111;
memory[4060]=8'b11111111;
memory[4061]=8'b11111111;
memory[4062]=8'b11111000;
memory[4063]=8'b00001111;
memory[4064]=8'b11111111;
memory[4065]=8'b11111000;
memory[4066]=8'b00000000;
memory[4067]=8'b11111111;
memory[4068]=8'b11111111;
memory[4069]=8'b11111111;
memory[4070]=8'b11111111;
memory[4071]=8'b11111111;
memory[4072]=8'b11111111;
memory[4073]=8'b11111111;
memory[4074]=8'b11111111;
memory[4075]=8'b11111111;
memory[4076]=8'b11111111;
memory[4077]=8'b11111111;
memory[4078]=8'b11111111;
memory[4079]=8'b11111111;
memory[4080]=8'b11111111;
memory[4081]=8'b11111111;
memory[4082]=8'b11111111;
memory[4083]=8'b11111111;
memory[4084]=8'b11111111;
memory[4085]=8'b11111111;
memory[4086]=8'b11111111;
memory[4087]=8'b11110000;
memory[4088]=8'b00000111;
memory[4089]=8'b11111111;
memory[4090]=8'b11111111;
memory[4091]=8'b11111100;
memory[4092]=8'b00000001;
memory[4093]=8'b11111111;
memory[4094]=8'b10000000;
memory[4095]=8'b01111111;
memory[4096]=8'b11111111;
memory[4097]=8'b11111111;
memory[4098]=8'b11111111;
memory[4099]=8'b11111111;
memory[4100]=8'b11111111;
memory[4101]=8'b11111111;
memory[4102]=8'b11110000;
memory[4103]=8'b00011111;
memory[4104]=8'b11111111;
memory[4105]=8'b11100000;
memory[4106]=8'b00000001;
memory[4107]=8'b11111111;
memory[4108]=8'b11111111;
memory[4109]=8'b00011111;
memory[4110]=8'b11111111;
memory[4111]=8'b11111111;
memory[4112]=8'b11111111;
memory[4113]=8'b11111111;
memory[4114]=8'b11111111;
memory[4115]=8'b11111111;
memory[4116]=8'b11111111;
memory[4117]=8'b11111111;
memory[4118]=8'b11111111;
memory[4119]=8'b11111111;
memory[4120]=8'b11111111;
memory[4121]=8'b11111111;
memory[4122]=8'b11111111;
memory[4123]=8'b11111111;
memory[4124]=8'b11111111;
memory[4125]=8'b11111111;
memory[4126]=8'b11111111;
memory[4127]=8'b11100000;
memory[4128]=8'b00011111;
memory[4129]=8'b11111111;
memory[4130]=8'b11111111;
memory[4131]=8'b11111111;
memory[4132]=8'b11000000;
memory[4133]=8'b00000000;
memory[4134]=8'b00000001;
memory[4135]=8'b11111111;
memory[4136]=8'b11111111;
memory[4137]=8'b11111111;
memory[4138]=8'b11111111;
memory[4139]=8'b11111111;
memory[4140]=8'b11111111;
memory[4141]=8'b11111111;
memory[4142]=8'b11110000;
memory[4143]=8'b00011111;
memory[4144]=8'b11111111;
memory[4145]=8'b10000000;
memory[4146]=8'b00000111;
memory[4147]=8'b11111111;
memory[4148]=8'b11111111;
memory[4149]=8'b11100011;
memory[4150]=8'b11111111;
memory[4151]=8'b11111111;
memory[4152]=8'b11111111;
memory[4153]=8'b11111111;
memory[4154]=8'b11111111;
memory[4155]=8'b11111111;
memory[4156]=8'b11111111;
memory[4157]=8'b11111111;
memory[4158]=8'b11111111;
memory[4159]=8'b11111111;
memory[4160]=8'b11111111;
memory[4161]=8'b11111111;
memory[4162]=8'b11111111;
memory[4163]=8'b11111111;
memory[4164]=8'b11111111;
memory[4165]=8'b11111111;
memory[4166]=8'b11111111;
memory[4167]=8'b11000000;
memory[4168]=8'b01111111;
memory[4169]=8'b11111111;
memory[4170]=8'b11111111;
memory[4171]=8'b11111111;
memory[4172]=8'b11111000;
memory[4173]=8'b01111110;
memory[4174]=8'b00000011;
memory[4175]=8'b11111111;
memory[4176]=8'b11111111;
memory[4177]=8'b11111111;
memory[4178]=8'b11111111;
memory[4179]=8'b11111111;
memory[4180]=8'b11111111;
memory[4181]=8'b11111111;
memory[4182]=8'b11100000;
memory[4183]=8'b00111111;
memory[4184]=8'b11111110;
memory[4185]=8'b00000000;
memory[4186]=8'b00011111;
memory[4187]=8'b11111111;
memory[4188]=8'b11111111;
memory[4189]=8'b11111000;
memory[4190]=8'b01111111;
memory[4191]=8'b11111111;
memory[4192]=8'b11111111;
memory[4193]=8'b11111111;
memory[4194]=8'b11111111;
memory[4195]=8'b11111111;
memory[4196]=8'b11111111;
memory[4197]=8'b11111111;
memory[4198]=8'b11111111;
memory[4199]=8'b11111111;
memory[4200]=8'b11111111;
memory[4201]=8'b11111111;
memory[4202]=8'b11111111;
memory[4203]=8'b11111111;
memory[4204]=8'b11111111;
memory[4205]=8'b11111111;
memory[4206]=8'b11111111;
memory[4207]=8'b11111101;
memory[4208]=8'b11111111;
memory[4209]=8'b11111111;
memory[4210]=8'b11111111;
memory[4211]=8'b11111111;
memory[4212]=8'b11111000;
memory[4213]=8'b00011111;
memory[4214]=8'b00000011;
memory[4215]=8'b11111111;
memory[4216]=8'b11111111;
memory[4217]=8'b11111111;
memory[4218]=8'b11111111;
memory[4219]=8'b11111111;
memory[4220]=8'b11111111;
memory[4221]=8'b11111111;
memory[4222]=8'b11000000;
memory[4223]=8'b01111111;
memory[4224]=8'b11111100;
memory[4225]=8'b00000000;
memory[4226]=8'b00111111;
memory[4227]=8'b11111111;
memory[4228]=8'b00111111;
memory[4229]=8'b11111111;
memory[4230]=8'b00011111;
memory[4231]=8'b11111111;
memory[4232]=8'b11111111;
memory[4233]=8'b11111111;
memory[4234]=8'b11111111;
memory[4235]=8'b11111111;
memory[4236]=8'b11111111;
memory[4237]=8'b11111111;
memory[4238]=8'b11111111;
memory[4239]=8'b11111111;
memory[4240]=8'b11111111;
memory[4241]=8'b11111111;
memory[4242]=8'b11111111;
memory[4243]=8'b11111111;
memory[4244]=8'b11111111;
memory[4245]=8'b11111111;
memory[4246]=8'b11111111;
memory[4247]=8'b11111111;
memory[4248]=8'b11111111;
memory[4249]=8'b11111111;
memory[4250]=8'b11111111;
memory[4251]=8'b11111111;
memory[4252]=8'b11111100;
memory[4253]=8'b00011111;
memory[4254]=8'b00000111;
memory[4255]=8'b11111111;
memory[4256]=8'b11111111;
memory[4257]=8'b11111111;
memory[4258]=8'b11111111;
memory[4259]=8'b11111111;
memory[4260]=8'b11111111;
memory[4261]=8'b11111111;
memory[4262]=8'b11000000;
memory[4263]=8'b01111111;
memory[4264]=8'b11111000;
memory[4265]=8'b00000000;
memory[4266]=8'b00111111;
memory[4267]=8'b11100111;
memory[4268]=8'b00111111;
memory[4269]=8'b11111111;
memory[4270]=8'b11100111;
memory[4271]=8'b11111111;
memory[4272]=8'b11111111;
memory[4273]=8'b11111111;
memory[4274]=8'b11111111;
memory[4275]=8'b11111111;
memory[4276]=8'b11111111;
memory[4277]=8'b11111111;
memory[4278]=8'b11111111;
memory[4279]=8'b11111111;
memory[4280]=8'b11111111;
memory[4281]=8'b11111111;
memory[4282]=8'b11111111;
memory[4283]=8'b11111111;
memory[4284]=8'b11111111;
memory[4285]=8'b11111111;
memory[4286]=8'b11111111;
memory[4287]=8'b11111111;
memory[4288]=8'b11111111;
memory[4289]=8'b11111111;
memory[4290]=8'b11111111;
memory[4291]=8'b11111111;
memory[4292]=8'b11111100;
memory[4293]=8'b00111111;
memory[4294]=8'b00001111;
memory[4295]=8'b11111111;
memory[4296]=8'b11111111;
memory[4297]=8'b11111111;
memory[4298]=8'b11111111;
memory[4299]=8'b11111111;
memory[4300]=8'b11111111;
memory[4301]=8'b11111111;
memory[4302]=8'b11000000;
memory[4303]=8'b01111111;
memory[4304]=8'b11110000;
memory[4305]=8'b00000000;
memory[4306]=8'b00001111;
memory[4307]=8'b11110000;
memory[4308]=8'b00111111;
memory[4309]=8'b11101111;
memory[4310]=8'b11111111;
memory[4311]=8'b11111111;
memory[4312]=8'b11111111;
memory[4313]=8'b11111111;
memory[4314]=8'b11111111;
memory[4315]=8'b11111111;
memory[4316]=8'b11111111;
memory[4317]=8'b11111111;
memory[4318]=8'b11111111;
memory[4319]=8'b11111111;
memory[4320]=8'b11111111;
memory[4321]=8'b11111111;
memory[4322]=8'b11111111;
memory[4323]=8'b11111111;
memory[4324]=8'b11111111;
memory[4325]=8'b11111111;
memory[4326]=8'b11111111;
memory[4327]=8'b11111111;
memory[4328]=8'b11111111;
memory[4329]=8'b11111111;
memory[4330]=8'b11111111;
memory[4331]=8'b11111111;
memory[4332]=8'b11111100;
memory[4333]=8'b00111110;
memory[4334]=8'b00001111;
memory[4335]=8'b11111111;
memory[4336]=8'b11111111;
memory[4337]=8'b11111111;
memory[4338]=8'b11111111;
memory[4339]=8'b11111111;
memory[4340]=8'b11111111;
memory[4341]=8'b11111111;
memory[4342]=8'b10000000;
memory[4343]=8'b01111111;
memory[4344]=8'b11110000;
memory[4345]=8'b00000000;
memory[4346]=8'b11111111;
memory[4347]=8'b11100000;
memory[4348]=8'b00111111;
memory[4349]=8'b11110011;
memory[4350]=8'b11111111;
memory[4351]=8'b11111111;
memory[4352]=8'b11111111;
memory[4353]=8'b11111111;
memory[4354]=8'b11111111;
memory[4355]=8'b11111111;
memory[4356]=8'b11111111;
memory[4357]=8'b11111111;
memory[4358]=8'b11111111;
memory[4359]=8'b11111111;
memory[4360]=8'b11111111;
memory[4361]=8'b11111111;
memory[4362]=8'b11111111;
memory[4363]=8'b11111111;
memory[4364]=8'b11111111;
memory[4365]=8'b11111111;
memory[4366]=8'b11111111;
memory[4367]=8'b11111111;
memory[4368]=8'b11111111;
memory[4369]=8'b11111111;
memory[4370]=8'b11111111;
memory[4371]=8'b11111111;
memory[4372]=8'b11111100;
memory[4373]=8'b00111110;
memory[4374]=8'b00001111;
memory[4375]=8'b11111111;
memory[4376]=8'b11111111;
memory[4377]=8'b11111111;
memory[4378]=8'b11111111;
memory[4379]=8'b11111111;
memory[4380]=8'b11111111;
memory[4381]=8'b11111111;
memory[4382]=8'b10000000;
memory[4383]=8'b11111111;
memory[4384]=8'b11100000;
memory[4385]=8'b00000000;
memory[4386]=8'b01111111;
memory[4387]=8'b11000000;
memory[4388]=8'b00000011;
memory[4389]=8'b11111001;
memory[4390]=8'b11011111;
memory[4391]=8'b11111111;
memory[4392]=8'b11111111;
memory[4393]=8'b11111111;
memory[4394]=8'b11111111;
memory[4395]=8'b11111111;
memory[4396]=8'b11111111;
memory[4397]=8'b11111111;
memory[4398]=8'b11111111;
memory[4399]=8'b11111111;
memory[4400]=8'b11111111;
memory[4401]=8'b11111111;
memory[4402]=8'b11111111;
memory[4403]=8'b11111111;
memory[4404]=8'b11111111;
memory[4405]=8'b11111111;
memory[4406]=8'b11111111;
memory[4407]=8'b11111111;
memory[4408]=8'b11111111;
memory[4409]=8'b11111111;
memory[4410]=8'b11111111;
memory[4411]=8'b11111111;
memory[4412]=8'b11111100;
memory[4413]=8'b00111110;
memory[4414]=8'b00011111;
memory[4415]=8'b11111111;
memory[4416]=8'b11111111;
memory[4417]=8'b11111111;
memory[4418]=8'b11111111;
memory[4419]=8'b11111111;
memory[4420]=8'b11111111;
memory[4421]=8'b11111111;
memory[4422]=8'b10000000;
memory[4423]=8'b11111111;
memory[4424]=8'b11000000;
memory[4425]=8'b00000000;
memory[4426]=8'b00011111;
memory[4427]=8'b10000000;
memory[4428]=8'b00000000;
memory[4429]=8'b01111001;
memory[4430]=8'b11001111;
memory[4431]=8'b10111111;
memory[4432]=8'b11111111;
memory[4433]=8'b11111111;
memory[4434]=8'b11111111;
memory[4435]=8'b11111111;
memory[4436]=8'b11111111;
memory[4437]=8'b11111111;
memory[4438]=8'b11111111;
memory[4439]=8'b11111111;
memory[4440]=8'b11111111;
memory[4441]=8'b11111111;
memory[4442]=8'b11111111;
memory[4443]=8'b11111111;
memory[4444]=8'b11111111;
memory[4445]=8'b11111111;
memory[4446]=8'b11111111;
memory[4447]=8'b11111111;
memory[4448]=8'b11111111;
memory[4449]=8'b11111111;
memory[4450]=8'b11111111;
memory[4451]=8'b11111111;
memory[4452]=8'b11111100;
memory[4453]=8'b00111100;
memory[4454]=8'b00011111;
memory[4455]=8'b11111111;
memory[4456]=8'b11111111;
memory[4457]=8'b11111111;
memory[4458]=8'b11111111;
memory[4459]=8'b11111111;
memory[4460]=8'b11111111;
memory[4461]=8'b11111111;
memory[4462]=8'b10000000;
memory[4463]=8'b01111111;
memory[4464]=8'b11000000;
memory[4465]=8'b00000000;
memory[4466]=8'b00001111;
memory[4467]=8'b10000000;
memory[4468]=8'b00000000;
memory[4469]=8'b00111100;
memory[4470]=8'b11001111;
memory[4471]=8'b10011111;
memory[4472]=8'b11111111;
memory[4473]=8'b11111111;
memory[4474]=8'b11111111;
memory[4475]=8'b11111111;
memory[4476]=8'b11111111;
memory[4477]=8'b11111111;
memory[4478]=8'b11111111;
memory[4479]=8'b11111111;
memory[4480]=8'b11111111;
memory[4481]=8'b11111111;
memory[4482]=8'b11111111;
memory[4483]=8'b11111111;
memory[4484]=8'b11111111;
memory[4485]=8'b11111111;
memory[4486]=8'b11111111;
memory[4487]=8'b11111111;
memory[4488]=8'b11111111;
memory[4489]=8'b11111111;
memory[4490]=8'b11111111;
memory[4491]=8'b11111111;
memory[4492]=8'b11111100;
memory[4493]=8'b01111100;
memory[4494]=8'b00011111;
memory[4495]=8'b11111111;
memory[4496]=8'b11111111;
memory[4497]=8'b11111111;
memory[4498]=8'b11111111;
memory[4499]=8'b11111111;
memory[4500]=8'b11111111;
memory[4501]=8'b11111111;
memory[4502]=8'b10000000;
memory[4503]=8'b01111111;
memory[4504]=8'b10000000;
memory[4505]=8'b00000000;
memory[4506]=8'b00001111;
memory[4507]=8'b11110000;
memory[4508]=8'b00000000;
memory[4509]=8'b00011100;
memory[4510]=8'b00001111;
memory[4511]=8'b00000111;
memory[4512]=8'b11111111;
memory[4513]=8'b11111111;
memory[4514]=8'b11111111;
memory[4515]=8'b11111111;
memory[4516]=8'b11111111;
memory[4517]=8'b11111111;
memory[4518]=8'b11111111;
memory[4519]=8'b11111111;
memory[4520]=8'b11111111;
memory[4521]=8'b11111111;
memory[4522]=8'b11111111;
memory[4523]=8'b11111111;
memory[4524]=8'b11111111;
memory[4525]=8'b11111111;
memory[4526]=8'b11111111;
memory[4527]=8'b11111111;
memory[4528]=8'b11111111;
memory[4529]=8'b11111111;
memory[4530]=8'b11111111;
memory[4531]=8'b11111111;
memory[4532]=8'b11111100;
memory[4533]=8'b01111100;
memory[4534]=8'b00011111;
memory[4535]=8'b11111111;
memory[4536]=8'b11111111;
memory[4537]=8'b11111111;
memory[4538]=8'b11111111;
memory[4539]=8'b11111111;
memory[4540]=8'b11111111;
memory[4541]=8'b11111111;
memory[4542]=8'b10000000;
memory[4543]=8'b00111111;
memory[4544]=8'b10000000;
memory[4545]=8'b00000000;
memory[4546]=8'b00001111;
memory[4547]=8'b11111110;
memory[4548]=8'b00000000;
memory[4549]=8'b00000000;
memory[4550]=8'b00000110;
memory[4551]=8'b00000011;
memory[4552]=8'b11111111;
memory[4553]=8'b11111111;
memory[4554]=8'b11111111;
memory[4555]=8'b11111111;
memory[4556]=8'b11111111;
memory[4557]=8'b11111111;
memory[4558]=8'b11111111;
memory[4559]=8'b11111111;
memory[4560]=8'b11111111;
memory[4561]=8'b11111111;
memory[4562]=8'b11111111;
memory[4563]=8'b11111111;
memory[4564]=8'b11111111;
memory[4565]=8'b11111111;
memory[4566]=8'b11111111;
memory[4567]=8'b11111111;
memory[4568]=8'b11111111;
memory[4569]=8'b11111111;
memory[4570]=8'b11111111;
memory[4571]=8'b11111111;
memory[4572]=8'b11111100;
memory[4573]=8'b01111100;
memory[4574]=8'b00111111;
memory[4575]=8'b11111111;
memory[4576]=8'b11111111;
memory[4577]=8'b11111111;
memory[4578]=8'b11111111;
memory[4579]=8'b11111111;
memory[4580]=8'b11111111;
memory[4581]=8'b11111111;
memory[4582]=8'b10000000;
memory[4583]=8'b00011110;
memory[4584]=8'b00000000;
memory[4585]=8'b00000000;
memory[4586]=8'b00000000;
memory[4587]=8'b00111111;
memory[4588]=8'b11111000;
memory[4589]=8'b00000000;
memory[4590]=8'b00000000;
memory[4591]=8'b00000000;
memory[4592]=8'b11111111;
memory[4593]=8'b11111111;
memory[4594]=8'b11111111;
memory[4595]=8'b11111111;
memory[4596]=8'b11111111;
memory[4597]=8'b11111111;
memory[4598]=8'b11111111;
memory[4599]=8'b11111111;
memory[4600]=8'b11111111;
memory[4601]=8'b11111111;
memory[4602]=8'b11111111;
memory[4603]=8'b11111111;
memory[4604]=8'b11111111;
memory[4605]=8'b11111111;
memory[4606]=8'b11111111;
memory[4607]=8'b11111111;
memory[4608]=8'b11111111;
memory[4609]=8'b11111111;
memory[4610]=8'b11111111;
memory[4611]=8'b11111111;
memory[4612]=8'b11111100;
memory[4613]=8'b01111100;
memory[4614]=8'b00111111;
memory[4615]=8'b11111111;
memory[4616]=8'b11111111;
memory[4617]=8'b11111111;
memory[4618]=8'b11111111;
memory[4619]=8'b11111111;
memory[4620]=8'b11111111;
memory[4621]=8'b11111111;
memory[4622]=8'b10000000;
memory[4623]=8'b00000000;
memory[4624]=8'b00000000;
memory[4625]=8'b00000000;
memory[4626]=8'b00000000;
memory[4627]=8'b00111111;
memory[4628]=8'b11111111;
memory[4629]=8'b10000000;
memory[4630]=8'b00000000;
memory[4631]=8'b00000000;
memory[4632]=8'b00111111;
memory[4633]=8'b11111111;
memory[4634]=8'b11111111;
memory[4635]=8'b11111111;
memory[4636]=8'b11111111;
memory[4637]=8'b11111111;
memory[4638]=8'b11111111;
memory[4639]=8'b11111111;
memory[4640]=8'b11111111;
memory[4641]=8'b11111111;
memory[4642]=8'b11111111;
memory[4643]=8'b11111111;
memory[4644]=8'b11111111;
memory[4645]=8'b11111111;
memory[4646]=8'b11111111;
memory[4647]=8'b11111111;
memory[4648]=8'b11111111;
memory[4649]=8'b11111111;
memory[4650]=8'b11111111;
memory[4651]=8'b11111111;
memory[4652]=8'b11111100;
memory[4653]=8'b01111000;
memory[4654]=8'b01111111;
memory[4655]=8'b11111111;
memory[4656]=8'b11111111;
memory[4657]=8'b11111111;
memory[4658]=8'b11111111;
memory[4659]=8'b11111111;
memory[4660]=8'b11111111;
memory[4661]=8'b11111111;
memory[4662]=8'b10000000;
memory[4663]=8'b00000000;
memory[4664]=8'b00000000;
memory[4665]=8'b00000000;
memory[4666]=8'b00000000;
memory[4667]=8'b11111111;
memory[4668]=8'b11111111;
memory[4669]=8'b11111111;
memory[4670]=8'b11111001;
memory[4671]=8'b11100000;
memory[4672]=8'b00001111;
memory[4673]=8'b11111111;
memory[4674]=8'b11111111;
memory[4675]=8'b11111111;
memory[4676]=8'b11111111;
memory[4677]=8'b11111111;
memory[4678]=8'b11111111;
memory[4679]=8'b11111111;
memory[4680]=8'b11111111;
memory[4681]=8'b11111111;
memory[4682]=8'b11111111;
memory[4683]=8'b11111111;
memory[4684]=8'b11111111;
memory[4685]=8'b11111111;
memory[4686]=8'b11111111;
memory[4687]=8'b11111111;
memory[4688]=8'b11111111;
memory[4689]=8'b11111111;
memory[4690]=8'b11111111;
memory[4691]=8'b11111111;
memory[4692]=8'b11111000;
memory[4693]=8'b01111000;
memory[4694]=8'b01111111;
memory[4695]=8'b11111111;
memory[4696]=8'b11111111;
memory[4697]=8'b11111111;
memory[4698]=8'b11111111;
memory[4699]=8'b11111111;
memory[4700]=8'b11111111;
memory[4701]=8'b11111111;
memory[4702]=8'b10000000;
memory[4703]=8'b00000000;
memory[4704]=8'b00000000;
memory[4705]=8'b00000000;
memory[4706]=8'b00000001;
memory[4707]=8'b11111100;
memory[4708]=8'b01111111;
memory[4709]=8'b11111111;
memory[4710]=8'b11111111;
memory[4711]=8'b11100000;
memory[4712]=8'b00000111;
memory[4713]=8'b11111111;
memory[4714]=8'b11111111;
memory[4715]=8'b11111111;
memory[4716]=8'b11111111;
memory[4717]=8'b11111111;
memory[4718]=8'b11111111;
memory[4719]=8'b11111111;
memory[4720]=8'b11111111;
memory[4721]=8'b11111111;
memory[4722]=8'b11111111;
memory[4723]=8'b11111111;
memory[4724]=8'b11111111;
memory[4725]=8'b11111111;
memory[4726]=8'b11111111;
memory[4727]=8'b11111111;
memory[4728]=8'b11111111;
memory[4729]=8'b11111111;
memory[4730]=8'b11111111;
memory[4731]=8'b11111111;
memory[4732]=8'b11111000;
memory[4733]=8'b11111000;
memory[4734]=8'b01111111;
memory[4735]=8'b11111111;
memory[4736]=8'b11111111;
memory[4737]=8'b11111111;
memory[4738]=8'b11111111;
memory[4739]=8'b11111111;
memory[4740]=8'b11111111;
memory[4741]=8'b11111111;
memory[4742]=8'b11000000;
memory[4743]=8'b00000000;
memory[4744]=8'b00000000;
memory[4745]=8'b00000000;
memory[4746]=8'b00000000;
memory[4747]=8'b00000000;
memory[4748]=8'b01111110;
memory[4749]=8'b00111111;
memory[4750]=8'b11111111;
memory[4751]=8'b11111000;
memory[4752]=8'b00000111;
memory[4753]=8'b11111111;
memory[4754]=8'b11111111;
memory[4755]=8'b11111111;
memory[4756]=8'b11111111;
memory[4757]=8'b11111111;
memory[4758]=8'b11111111;
memory[4759]=8'b11111111;
memory[4760]=8'b11111111;
memory[4761]=8'b11111111;
memory[4762]=8'b11111111;
memory[4763]=8'b11111111;
memory[4764]=8'b11111111;
memory[4765]=8'b11111111;
memory[4766]=8'b11111111;
memory[4767]=8'b11111111;
memory[4768]=8'b11111111;
memory[4769]=8'b11111111;
memory[4770]=8'b11111111;
memory[4771]=8'b11111111;
memory[4772]=8'b11111000;
memory[4773]=8'b11111000;
memory[4774]=8'b11111111;
memory[4775]=8'b11111111;
memory[4776]=8'b11111111;
memory[4777]=8'b11111111;
memory[4778]=8'b11111111;
memory[4779]=8'b11111111;
memory[4780]=8'b11111111;
memory[4781]=8'b11111111;
memory[4782]=8'b11100000;
memory[4783]=8'b00000000;
memory[4784]=8'b00000000;
memory[4785]=8'b00000000;
memory[4786]=8'b00000000;
memory[4787]=8'b00000000;
memory[4788]=8'b00000000;
memory[4789]=8'b00011111;
memory[4790]=8'b11110000;
memory[4791]=8'b11111110;
memory[4792]=8'b00000111;
memory[4793]=8'b11111111;
memory[4794]=8'b11111111;
memory[4795]=8'b11111111;
memory[4796]=8'b11111111;
memory[4797]=8'b11111111;
memory[4798]=8'b11111111;
memory[4799]=8'b11111111;
memory[4800]=8'b11111111;
memory[4801]=8'b11111111;
memory[4802]=8'b11111111;
memory[4803]=8'b11111111;
memory[4804]=8'b11111111;
memory[4805]=8'b11111111;
memory[4806]=8'b11111111;
memory[4807]=8'b11111111;
memory[4808]=8'b11111111;
memory[4809]=8'b11111111;
memory[4810]=8'b11111111;
memory[4811]=8'b11111111;
memory[4812]=8'b11111000;
memory[4813]=8'b11110000;
memory[4814]=8'b11111111;
memory[4815]=8'b11111111;
memory[4816]=8'b11111111;
memory[4817]=8'b11111111;
memory[4818]=8'b11111111;
memory[4819]=8'b11111111;
memory[4820]=8'b11111111;
memory[4821]=8'b11111111;
memory[4822]=8'b11111000;
memory[4823]=8'b00000000;
memory[4824]=8'b00000000;
memory[4825]=8'b00001111;
memory[4826]=8'b11000000;
memory[4827]=8'b00000000;
memory[4828]=8'b00000000;
memory[4829]=8'b00000000;
memory[4830]=8'b00000000;
memory[4831]=8'b00011111;
memory[4832]=8'b11000011;
memory[4833]=8'b11111111;
memory[4834]=8'b11111111;
memory[4835]=8'b11111111;
memory[4836]=8'b11111111;
memory[4837]=8'b11111111;
memory[4838]=8'b11111111;
memory[4839]=8'b11111111;
memory[4840]=8'b11111111;
memory[4841]=8'b11111111;
memory[4842]=8'b11111111;
memory[4843]=8'b11111111;
memory[4844]=8'b11111111;
memory[4845]=8'b11111111;
memory[4846]=8'b11111111;
memory[4847]=8'b11111111;
memory[4848]=8'b11111111;
memory[4849]=8'b11111111;
memory[4850]=8'b11111111;
memory[4851]=8'b11111111;
memory[4852]=8'b11111000;
memory[4853]=8'b11110000;
memory[4854]=8'b11111111;
memory[4855]=8'b11111111;
memory[4856]=8'b11111111;
memory[4857]=8'b11111111;
memory[4858]=8'b11111111;
memory[4859]=8'b11111111;
memory[4860]=8'b11111111;
memory[4861]=8'b11111111;
memory[4862]=8'b11111110;
memory[4863]=8'b00000000;
memory[4864]=8'b00000001;
memory[4865]=8'b11111111;
memory[4866]=8'b11111100;
memory[4867]=8'b00000000;
memory[4868]=8'b00000000;
memory[4869]=8'b00000011;
memory[4870]=8'b11111111;
memory[4871]=8'b00000011;
memory[4872]=8'b11111001;
memory[4873]=8'b11111111;
memory[4874]=8'b11111111;
memory[4875]=8'b11111111;
memory[4876]=8'b11111111;
memory[4877]=8'b11111111;
memory[4878]=8'b11111111;
memory[4879]=8'b11111111;
memory[4880]=8'b11111111;
memory[4881]=8'b11111111;
memory[4882]=8'b11111111;
memory[4883]=8'b11111111;
memory[4884]=8'b11111111;
memory[4885]=8'b11111111;
memory[4886]=8'b11111111;
memory[4887]=8'b11111111;
memory[4888]=8'b11111111;
memory[4889]=8'b11111111;
memory[4890]=8'b11111111;
memory[4891]=8'b11111111;
memory[4892]=8'b11110001;
memory[4893]=8'b11110000;
memory[4894]=8'b11111111;
memory[4895]=8'b11111111;
memory[4896]=8'b11111111;
memory[4897]=8'b11111111;
memory[4898]=8'b11111111;
memory[4899]=8'b11111111;
memory[4900]=8'b11111111;
memory[4901]=8'b11111111;
memory[4902]=8'b11111111;
memory[4903]=8'b11100000;
memory[4904]=8'b00011111;
memory[4905]=8'b11110000;
memory[4906]=8'b00111111;
memory[4907]=8'b11000000;
memory[4908]=8'b00000000;
memory[4909]=8'b00111111;
memory[4910]=8'b11111111;
memory[4911]=8'b11000000;
memory[4912]=8'b01111111;
memory[4913]=8'b11111111;
memory[4914]=8'b11111111;
memory[4915]=8'b11111111;
memory[4916]=8'b11111111;
memory[4917]=8'b11111111;
memory[4918]=8'b11111111;
memory[4919]=8'b11111111;
memory[4920]=8'b11111111;
memory[4921]=8'b11111111;
memory[4922]=8'b11111111;
memory[4923]=8'b11111111;
memory[4924]=8'b11111111;
memory[4925]=8'b11111111;
memory[4926]=8'b11111111;
memory[4927]=8'b11111111;
memory[4928]=8'b11111111;
memory[4929]=8'b11111111;
memory[4930]=8'b11111111;
memory[4931]=8'b11111111;
memory[4932]=8'b11110001;
memory[4933]=8'b11110000;
memory[4934]=8'b11111111;
memory[4935]=8'b11111111;
memory[4936]=8'b11111111;
memory[4937]=8'b11111111;
memory[4938]=8'b11111111;
memory[4939]=8'b11111111;
memory[4940]=8'b11111111;
memory[4941]=8'b11111111;
memory[4942]=8'b11111111;
memory[4943]=8'b11111111;
memory[4944]=8'b11111110;
memory[4945]=8'b00000110;
memory[4946]=8'b00000011;
memory[4947]=8'b11111110;
memory[4948]=8'b00111111;
memory[4949]=8'b11111100;
memory[4950]=8'b00000111;
memory[4951]=8'b11110000;
memory[4952]=8'b00011111;
memory[4953]=8'b11111111;
memory[4954]=8'b11111111;
memory[4955]=8'b11111111;
memory[4956]=8'b11111111;
memory[4957]=8'b11111111;
memory[4958]=8'b11111111;
memory[4959]=8'b11111111;
memory[4960]=8'b11111111;
memory[4961]=8'b11111111;
memory[4962]=8'b11111111;
memory[4963]=8'b11111111;
memory[4964]=8'b11111111;
memory[4965]=8'b11111111;
memory[4966]=8'b11111111;
memory[4967]=8'b11111111;
memory[4968]=8'b11111111;
memory[4969]=8'b11111111;
memory[4970]=8'b11111111;
memory[4971]=8'b11111111;
memory[4972]=8'b11110001;
memory[4973]=8'b11100000;
memory[4974]=8'b11111111;
memory[4975]=8'b11111111;
memory[4976]=8'b11111111;
memory[4977]=8'b11111111;
memory[4978]=8'b11111111;
memory[4979]=8'b11111111;
memory[4980]=8'b11111111;
memory[4981]=8'b11111111;
memory[4982]=8'b11111111;
memory[4983]=8'b11111111;
memory[4984]=8'b11111111;
memory[4985]=8'b11111111;
memory[4986]=8'b11111000;
memory[4987]=8'b01111111;
memory[4988]=8'b11111111;
memory[4989]=8'b11001111;
memory[4990]=8'b11111111;
memory[4991]=8'b11111000;
memory[4992]=8'b00001111;
memory[4993]=8'b11111111;
memory[4994]=8'b11111111;
memory[4995]=8'b11111111;
memory[4996]=8'b11111111;
memory[4997]=8'b11111111;
memory[4998]=8'b11111111;
memory[4999]=8'b11111111;
memory[5000]=8'b11111111;
memory[5001]=8'b11111111;
memory[5002]=8'b11111111;
memory[5003]=8'b11111111;
memory[5004]=8'b11111111;
memory[5005]=8'b11111111;
memory[5006]=8'b11111111;
memory[5007]=8'b11111111;
memory[5008]=8'b11111111;
memory[5009]=8'b11111111;
memory[5010]=8'b11111111;
memory[5011]=8'b11111111;
memory[5012]=8'b11110001;
memory[5013]=8'b11100000;
memory[5014]=8'b11111111;
memory[5015]=8'b11111111;
memory[5016]=8'b11111111;
memory[5017]=8'b11111111;
memory[5018]=8'b11111111;
memory[5019]=8'b11111111;
memory[5020]=8'b11111111;
memory[5021]=8'b11111111;
memory[5022]=8'b11111111;
memory[5023]=8'b11111111;
memory[5024]=8'b11111111;
memory[5025]=8'b11111111;
memory[5026]=8'b11111110;
memory[5027]=8'b00000000;
memory[5028]=8'b00000000;
memory[5029]=8'b01111111;
memory[5030]=8'b11111111;
memory[5031]=8'b11111110;
memory[5032]=8'b00000111;
memory[5033]=8'b11111111;
memory[5034]=8'b11111111;
memory[5035]=8'b11111111;
memory[5036]=8'b11111111;
memory[5037]=8'b11111111;
memory[5038]=8'b11111111;
memory[5039]=8'b11111111;
memory[5040]=8'b11111111;
memory[5041]=8'b11111111;
memory[5042]=8'b11111111;
memory[5043]=8'b11111111;
memory[5044]=8'b11111111;
memory[5045]=8'b11111111;
memory[5046]=8'b11111111;
memory[5047]=8'b11111111;
memory[5048]=8'b11111111;
memory[5049]=8'b11111111;
memory[5050]=8'b11111111;
memory[5051]=8'b11111111;
memory[5052]=8'b11110001;
memory[5053]=8'b11100001;
memory[5054]=8'b11111111;
memory[5055]=8'b11111111;
memory[5056]=8'b11111111;
memory[5057]=8'b11111111;
memory[5058]=8'b11111111;
memory[5059]=8'b11111111;
memory[5060]=8'b11111111;
memory[5061]=8'b11111111;
memory[5062]=8'b11111111;
memory[5063]=8'b11111111;
memory[5064]=8'b11111111;
memory[5065]=8'b11111111;
memory[5066]=8'b11111111;
memory[5067]=8'b10000011;
memory[5068]=8'b10000111;
memory[5069]=8'b11111111;
memory[5070]=8'b11111111;
memory[5071]=8'b11111111;
memory[5072]=8'b10000011;
memory[5073]=8'b11111111;
memory[5074]=8'b11111111;
memory[5075]=8'b11111111;
memory[5076]=8'b11111111;
memory[5077]=8'b11111111;
memory[5078]=8'b11111111;
memory[5079]=8'b11111111;
memory[5080]=8'b11111111;
memory[5081]=8'b11111111;
memory[5082]=8'b11111111;
memory[5083]=8'b11111111;
memory[5084]=8'b11111111;
memory[5085]=8'b11111111;
memory[5086]=8'b11111111;
memory[5087]=8'b11111111;
memory[5088]=8'b11111111;
memory[5089]=8'b11111111;
memory[5090]=8'b11111111;
memory[5091]=8'b11111111;
memory[5092]=8'b11110011;
memory[5093]=8'b11100001;
memory[5094]=8'b11111111;
memory[5095]=8'b11111111;
memory[5096]=8'b11111111;
memory[5097]=8'b11111111;
memory[5098]=8'b11111111;
memory[5099]=8'b11111111;
memory[5100]=8'b11111111;
memory[5101]=8'b11111111;
memory[5102]=8'b11111111;
memory[5103]=8'b11111111;
memory[5104]=8'b11111111;
memory[5105]=8'b11111111;
memory[5106]=8'b11111111;
memory[5107]=8'b10000111;
memory[5108]=8'b10000111;
memory[5109]=8'b11111111;
memory[5110]=8'b11111111;
memory[5111]=8'b11111111;
memory[5112]=8'b11111111;
memory[5113]=8'b11111111;
memory[5114]=8'b11111111;
memory[5115]=8'b11111111;
memory[5116]=8'b11111111;
memory[5117]=8'b11111111;
memory[5118]=8'b11111111;
memory[5119]=8'b11111111;
memory[5120]=8'b11111111;
memory[5121]=8'b11111111;
memory[5122]=8'b11111111;
memory[5123]=8'b11111111;
memory[5124]=8'b11111111;
memory[5125]=8'b11111111;
memory[5126]=8'b11111111;
memory[5127]=8'b11111111;
memory[5128]=8'b11111111;
memory[5129]=8'b11111111;
memory[5130]=8'b11111111;
memory[5131]=8'b11111111;
memory[5132]=8'b11100011;
memory[5133]=8'b11100001;
memory[5134]=8'b11111111;
memory[5135]=8'b11111111;
memory[5136]=8'b11111111;
memory[5137]=8'b11111111;
memory[5138]=8'b11111111;
memory[5139]=8'b11111111;
memory[5140]=8'b11111111;
memory[5141]=8'b11111111;
memory[5142]=8'b11111111;
memory[5143]=8'b11111111;
memory[5144]=8'b11111111;
memory[5145]=8'b11111111;
memory[5146]=8'b11111111;
memory[5147]=8'b11000111;
memory[5148]=8'b10000111;
memory[5149]=8'b11111111;
memory[5150]=8'b11111111;
memory[5151]=8'b11111111;
memory[5152]=8'b11111111;
memory[5153]=8'b11111111;
memory[5154]=8'b11111111;
memory[5155]=8'b11111111;
memory[5156]=8'b11111111;
memory[5157]=8'b11111111;
memory[5158]=8'b11111111;
memory[5159]=8'b11111111;
memory[5160]=8'b11111111;
memory[5161]=8'b11111111;
memory[5162]=8'b11111111;
memory[5163]=8'b11111111;
memory[5164]=8'b11111111;
memory[5165]=8'b11111111;
memory[5166]=8'b11111111;
memory[5167]=8'b11111111;
memory[5168]=8'b11111111;
memory[5169]=8'b11111111;
memory[5170]=8'b11111111;
memory[5171]=8'b11111111;
memory[5172]=8'b11100011;
memory[5173]=8'b11000011;
memory[5174]=8'b11111111;
memory[5175]=8'b11111111;
memory[5176]=8'b11111111;
memory[5177]=8'b11111111;
memory[5178]=8'b11111111;
memory[5179]=8'b11111111;
memory[5180]=8'b11111111;
memory[5181]=8'b11111111;
memory[5182]=8'b11111111;
memory[5183]=8'b11111111;
memory[5184]=8'b11111111;
memory[5185]=8'b11111111;
memory[5186]=8'b11111111;
memory[5187]=8'b11000111;
memory[5188]=8'b11000111;
memory[5189]=8'b11111111;
memory[5190]=8'b11111111;
memory[5191]=8'b11111111;
memory[5192]=8'b11111111;
memory[5193]=8'b11111111;
memory[5194]=8'b11111111;
memory[5195]=8'b11111111;
memory[5196]=8'b11111111;
memory[5197]=8'b11111111;
memory[5198]=8'b11111111;
memory[5199]=8'b11111111;
memory[5200]=8'b11111111;
memory[5201]=8'b11111111;
memory[5202]=8'b11111111;
memory[5203]=8'b11111111;
memory[5204]=8'b11111111;
memory[5205]=8'b11111111;
memory[5206]=8'b11111111;
memory[5207]=8'b11111111;
memory[5208]=8'b11111111;
memory[5209]=8'b11111111;
memory[5210]=8'b11111111;
memory[5211]=8'b11111111;
memory[5212]=8'b11100011;
memory[5213]=8'b11000011;
memory[5214]=8'b11111111;
memory[5215]=8'b11111111;
memory[5216]=8'b11111111;
memory[5217]=8'b11111111;
memory[5218]=8'b11111111;
memory[5219]=8'b11111111;
memory[5220]=8'b11111111;
memory[5221]=8'b11111111;
memory[5222]=8'b11111111;
memory[5223]=8'b11111111;
memory[5224]=8'b11111111;
memory[5225]=8'b11111111;
memory[5226]=8'b11111111;
memory[5227]=8'b11000011;
memory[5228]=8'b11000111;
memory[5229]=8'b11111111;
memory[5230]=8'b11111111;
memory[5231]=8'b11111111;
memory[5232]=8'b11111111;
memory[5233]=8'b11111111;
memory[5234]=8'b11111111;
memory[5235]=8'b11111111;
memory[5236]=8'b11111111;
memory[5237]=8'b11111111;
memory[5238]=8'b11111111;
memory[5239]=8'b11111111;
memory[5240]=8'b11111111;
memory[5241]=8'b11111111;
memory[5242]=8'b11111111;
memory[5243]=8'b11111111;
memory[5244]=8'b11111111;
memory[5245]=8'b11111111;
memory[5246]=8'b11111111;
memory[5247]=8'b11111111;
memory[5248]=8'b11111111;
memory[5249]=8'b11111111;
memory[5250]=8'b11111111;
memory[5251]=8'b11111111;
memory[5252]=8'b11100011;
memory[5253]=8'b10000111;
memory[5254]=8'b11111111;
memory[5255]=8'b11111111;
memory[5256]=8'b11111111;
memory[5257]=8'b11111111;
memory[5258]=8'b11111111;
memory[5259]=8'b11111111;
memory[5260]=8'b11111111;
memory[5261]=8'b11111111;
memory[5262]=8'b11111111;
memory[5263]=8'b11111111;
memory[5264]=8'b11111111;
memory[5265]=8'b11111111;
memory[5266]=8'b11111111;
memory[5267]=8'b11100011;
memory[5268]=8'b11000111;
memory[5269]=8'b11111111;
memory[5270]=8'b11111111;
memory[5271]=8'b11111111;
memory[5272]=8'b11111111;
memory[5273]=8'b11111111;
memory[5274]=8'b11111111;
memory[5275]=8'b11111111;
memory[5276]=8'b11111111;
memory[5277]=8'b11111111;
memory[5278]=8'b11111111;
memory[5279]=8'b11111111;
memory[5280]=8'b11111111;
memory[5281]=8'b11111111;
memory[5282]=8'b11111111;
memory[5283]=8'b11111111;
memory[5284]=8'b11111111;
memory[5285]=8'b11111111;
memory[5286]=8'b11111111;
memory[5287]=8'b11111111;
memory[5288]=8'b11111111;
memory[5289]=8'b11111111;
memory[5290]=8'b11111111;
memory[5291]=8'b11111111;
memory[5292]=8'b11100011;
memory[5293]=8'b10000111;
memory[5294]=8'b11111111;
memory[5295]=8'b11111111;
memory[5296]=8'b11111111;
memory[5297]=8'b11111111;
memory[5298]=8'b11111111;
memory[5299]=8'b11111111;
memory[5300]=8'b11111111;
memory[5301]=8'b11111111;
memory[5302]=8'b11111111;
memory[5303]=8'b11111111;
memory[5304]=8'b11111111;
memory[5305]=8'b11111111;
memory[5306]=8'b11111111;
memory[5307]=8'b11100011;
memory[5308]=8'b11000111;
memory[5309]=8'b11111111;
memory[5310]=8'b11111111;
memory[5311]=8'b11111111;
memory[5312]=8'b11111111;
memory[5313]=8'b11111111;
memory[5314]=8'b11111111;
memory[5315]=8'b11111111;
memory[5316]=8'b11111111;
memory[5317]=8'b11111111;
memory[5318]=8'b11111111;
memory[5319]=8'b11111111;
memory[5320]=8'b11111111;
memory[5321]=8'b11111111;
memory[5322]=8'b11111111;
memory[5323]=8'b11111111;
memory[5324]=8'b11111111;
memory[5325]=8'b11111111;
memory[5326]=8'b11111111;
memory[5327]=8'b11111111;
memory[5328]=8'b11111111;
memory[5329]=8'b11111111;
memory[5330]=8'b11111111;
memory[5331]=8'b11111111;
memory[5332]=8'b11000011;
memory[5333]=8'b10000111;
memory[5334]=8'b11111111;
memory[5335]=8'b11111111;
memory[5336]=8'b11111111;
memory[5337]=8'b11111111;
memory[5338]=8'b11111111;
memory[5339]=8'b11111111;
memory[5340]=8'b11111111;
memory[5341]=8'b11111111;
memory[5342]=8'b11111111;
memory[5343]=8'b11111111;
memory[5344]=8'b11111111;
memory[5345]=8'b11111111;
memory[5346]=8'b11111111;
memory[5347]=8'b11100001;
memory[5348]=8'b11000111;
memory[5349]=8'b11111111;
memory[5350]=8'b11111111;
memory[5351]=8'b11111111;
memory[5352]=8'b11111111;
memory[5353]=8'b11111111;
memory[5354]=8'b11111111;
memory[5355]=8'b11111111;
memory[5356]=8'b11111111;
memory[5357]=8'b11111111;
memory[5358]=8'b11111111;
memory[5359]=8'b11111111;
memory[5360]=8'b11111111;
memory[5361]=8'b11111111;
memory[5362]=8'b11111111;
memory[5363]=8'b11111111;
memory[5364]=8'b11111111;
memory[5365]=8'b11111111;
memory[5366]=8'b11111111;
memory[5367]=8'b11111111;
memory[5368]=8'b11111111;
memory[5369]=8'b11111111;
memory[5370]=8'b11111111;
memory[5371]=8'b11111111;
memory[5372]=8'b11000111;
memory[5373]=8'b10000011;
memory[5374]=8'b11111111;
memory[5375]=8'b11111111;
memory[5376]=8'b11111111;
memory[5377]=8'b11111111;
memory[5378]=8'b11111111;
memory[5379]=8'b11111111;
memory[5380]=8'b11111111;
memory[5381]=8'b11111111;
memory[5382]=8'b11111111;
memory[5383]=8'b11111111;
memory[5384]=8'b11111111;
memory[5385]=8'b11111111;
memory[5386]=8'b11111111;
memory[5387]=8'b11110001;
memory[5388]=8'b11100111;
memory[5389]=8'b11111111;
memory[5390]=8'b11111111;
memory[5391]=8'b11111111;
memory[5392]=8'b11111111;
memory[5393]=8'b11111111;
memory[5394]=8'b11111111;
memory[5395]=8'b11111111;
memory[5396]=8'b11111111;
memory[5397]=8'b11111111;
memory[5398]=8'b11111111;
memory[5399]=8'b11111111;
memory[5400]=8'b11111111;
memory[5401]=8'b11111111;
memory[5402]=8'b11111111;
memory[5403]=8'b11111111;
memory[5404]=8'b11111111;
memory[5405]=8'b11111111;
memory[5406]=8'b11111111;
memory[5407]=8'b11111111;
memory[5408]=8'b11111111;
memory[5409]=8'b11111111;
memory[5410]=8'b11111111;
memory[5411]=8'b11111111;
memory[5412]=8'b11000011;
memory[5413]=8'b10000011;
memory[5414]=8'b11111111;
memory[5415]=8'b11111111;
memory[5416]=8'b11111111;
memory[5417]=8'b11111111;
memory[5418]=8'b11111111;
memory[5419]=8'b11111111;
memory[5420]=8'b11111111;
memory[5421]=8'b11111111;
memory[5422]=8'b11111111;
memory[5423]=8'b11111111;
memory[5424]=8'b11111111;
memory[5425]=8'b11111111;
memory[5426]=8'b11111111;
memory[5427]=8'b11110001;
memory[5428]=8'b11100111;
memory[5429]=8'b11111111;
memory[5430]=8'b11111111;
memory[5431]=8'b11111111;
memory[5432]=8'b11111111;
memory[5433]=8'b11111111;
memory[5434]=8'b11111111;
memory[5435]=8'b11111111;
memory[5436]=8'b11111111;
memory[5437]=8'b11111111;
memory[5438]=8'b11111111;
memory[5439]=8'b11111111;
memory[5440]=8'b11111111;
memory[5441]=8'b11111111;
memory[5442]=8'b11111111;
memory[5443]=8'b11111111;
memory[5444]=8'b11111111;
memory[5445]=8'b11111111;
memory[5446]=8'b11111111;
memory[5447]=8'b11111111;
memory[5448]=8'b11111111;
memory[5449]=8'b11111111;
memory[5450]=8'b11111111;
memory[5451]=8'b11111111;
memory[5452]=8'b11000011;
memory[5453]=8'b10000011;
memory[5454]=8'b11111111;
memory[5455]=8'b11111111;
memory[5456]=8'b11111111;
memory[5457]=8'b11111111;
memory[5458]=8'b11111111;
memory[5459]=8'b11111111;
memory[5460]=8'b11111111;
memory[5461]=8'b11111111;
memory[5462]=8'b11111111;
memory[5463]=8'b11111111;
memory[5464]=8'b11111111;
memory[5465]=8'b11111111;
memory[5466]=8'b11111111;
memory[5467]=8'b11110001;
memory[5468]=8'b11100111;
memory[5469]=8'b11111111;
memory[5470]=8'b11111111;
memory[5471]=8'b11111111;
memory[5472]=8'b11111111;
memory[5473]=8'b11111111;
memory[5474]=8'b11111111;
memory[5475]=8'b11111111;
memory[5476]=8'b11111111;
memory[5477]=8'b11111111;
memory[5478]=8'b11111111;
memory[5479]=8'b11111111;
memory[5480]=8'b11111111;
memory[5481]=8'b11111111;
memory[5482]=8'b11111111;
memory[5483]=8'b11111111;
memory[5484]=8'b11111111;
memory[5485]=8'b11111111;
memory[5486]=8'b11111111;
memory[5487]=8'b11111111;
memory[5488]=8'b11111111;
memory[5489]=8'b11111111;
memory[5490]=8'b11111111;
memory[5491]=8'b11111111;
memory[5492]=8'b10000011;
memory[5493]=8'b10000011;
memory[5494]=8'b11111111;
memory[5495]=8'b11111111;
memory[5496]=8'b11111111;
memory[5497]=8'b11111111;
memory[5498]=8'b11111111;
memory[5499]=8'b11111111;
memory[5500]=8'b11111111;
memory[5501]=8'b11111111;
memory[5502]=8'b11111111;
memory[5503]=8'b11111111;
memory[5504]=8'b11111111;
memory[5505]=8'b11111111;
memory[5506]=8'b11111111;
memory[5507]=8'b11111001;
memory[5508]=8'b11100111;
memory[5509]=8'b11111111;
memory[5510]=8'b11111111;
memory[5511]=8'b11111111;
memory[5512]=8'b11111111;
memory[5513]=8'b11111111;
memory[5514]=8'b11111111;
memory[5515]=8'b11111111;
memory[5516]=8'b11111111;
memory[5517]=8'b11111111;
memory[5518]=8'b11111111;
memory[5519]=8'b11111111;
memory[5520]=8'b11111111;
memory[5521]=8'b11111111;
memory[5522]=8'b11111111;
memory[5523]=8'b11111111;
memory[5524]=8'b11111111;
memory[5525]=8'b11111111;
memory[5526]=8'b11111111;
memory[5527]=8'b11111111;
memory[5528]=8'b11111111;
memory[5529]=8'b11111111;
memory[5530]=8'b11111111;
memory[5531]=8'b11111111;
memory[5532]=8'b10000001;
memory[5533]=8'b10000001;
memory[5534]=8'b11111111;
memory[5535]=8'b11111111;
memory[5536]=8'b11111111;
memory[5537]=8'b11111111;
memory[5538]=8'b11111111;
memory[5539]=8'b11111111;
memory[5540]=8'b11111111;
memory[5541]=8'b11111111;
memory[5542]=8'b11111111;
memory[5543]=8'b11111111;
memory[5544]=8'b11111111;
memory[5545]=8'b11111111;
memory[5546]=8'b11111111;
memory[5547]=8'b11111000;
memory[5548]=8'b11100011;
memory[5549]=8'b11111111;
memory[5550]=8'b11111111;
memory[5551]=8'b11111111;
memory[5552]=8'b11111111;
memory[5553]=8'b11111111;
memory[5554]=8'b11111111;
memory[5555]=8'b11111111;
memory[5556]=8'b11111111;
memory[5557]=8'b11111111;
memory[5558]=8'b11111111;
memory[5559]=8'b11111111;
memory[5560]=8'b11111111;
memory[5561]=8'b11111111;
memory[5562]=8'b11111111;
memory[5563]=8'b11111111;
memory[5564]=8'b11111111;
memory[5565]=8'b11111111;
memory[5566]=8'b11111111;
memory[5567]=8'b11111111;
memory[5568]=8'b11111111;
memory[5569]=8'b11111111;
memory[5570]=8'b11111111;
memory[5571]=8'b11111111;
memory[5572]=8'b10000000;
memory[5573]=8'b10000001;
memory[5574]=8'b11111111;
memory[5575]=8'b11111111;
memory[5576]=8'b11111111;
memory[5577]=8'b11111111;
memory[5578]=8'b11111111;
memory[5579]=8'b11111111;
memory[5580]=8'b11111111;
memory[5581]=8'b11111111;
memory[5582]=8'b11111111;
memory[5583]=8'b11111111;
memory[5584]=8'b11111111;
memory[5585]=8'b11111111;
memory[5586]=8'b11111111;
memory[5587]=8'b11111000;
memory[5588]=8'b11110011;
memory[5589]=8'b11111111;
memory[5590]=8'b11111111;
memory[5591]=8'b11111111;
memory[5592]=8'b11111111;
memory[5593]=8'b11111111;
memory[5594]=8'b11111111;
memory[5595]=8'b11111111;
memory[5596]=8'b11111111;
memory[5597]=8'b11111111;
memory[5598]=8'b11111111;
memory[5599]=8'b11111111;
memory[5600]=8'b11111111;
memory[5601]=8'b11111111;
memory[5602]=8'b11111111;
memory[5603]=8'b11111111;
memory[5604]=8'b11111111;
memory[5605]=8'b11111111;
memory[5606]=8'b11111111;
memory[5607]=8'b11111111;
memory[5608]=8'b11111111;
memory[5609]=8'b11111111;
memory[5610]=8'b11111111;
memory[5611]=8'b11111111;
memory[5612]=8'b11000000;
memory[5613]=8'b11000011;
memory[5614]=8'b11111111;
memory[5615]=8'b11111111;
memory[5616]=8'b11111111;
memory[5617]=8'b11111111;
memory[5618]=8'b11111111;
memory[5619]=8'b11111111;
memory[5620]=8'b11111111;
memory[5621]=8'b11111111;
memory[5622]=8'b11111111;
memory[5623]=8'b11111111;
memory[5624]=8'b11111111;
memory[5625]=8'b11111111;
memory[5626]=8'b11111111;
memory[5627]=8'b11111000;
memory[5628]=8'b11110011;
memory[5629]=8'b11111111;
memory[5630]=8'b11111111;
memory[5631]=8'b11111111;
memory[5632]=8'b11111111;
memory[5633]=8'b11111111;
memory[5634]=8'b11111111;
memory[5635]=8'b11111111;
memory[5636]=8'b11111111;
memory[5637]=8'b11111111;
memory[5638]=8'b11111111;
memory[5639]=8'b11111111;
memory[5640]=8'b11111111;
memory[5641]=8'b11111111;
memory[5642]=8'b11111111;
memory[5643]=8'b11111111;
memory[5644]=8'b11111111;
memory[5645]=8'b11111111;
memory[5646]=8'b11111111;
memory[5647]=8'b11111111;
memory[5648]=8'b11111111;
memory[5649]=8'b11111111;
memory[5650]=8'b11111111;
memory[5651]=8'b11111111;
memory[5652]=8'b11000000;
memory[5653]=8'b11000011;
memory[5654]=8'b11111111;
memory[5655]=8'b11111111;
memory[5656]=8'b11111111;
memory[5657]=8'b11111111;
memory[5658]=8'b11111111;
memory[5659]=8'b11111111;
memory[5660]=8'b11111111;
memory[5661]=8'b11111111;
memory[5662]=8'b11111111;
memory[5663]=8'b11111111;
memory[5664]=8'b11111111;
memory[5665]=8'b11111111;
memory[5666]=8'b11111111;
memory[5667]=8'b11111000;
memory[5668]=8'b11110011;
memory[5669]=8'b11111111;
memory[5670]=8'b11111111;
memory[5671]=8'b11111111;
memory[5672]=8'b11111111;
memory[5673]=8'b11111111;
memory[5674]=8'b11111111;
memory[5675]=8'b11111111;
memory[5676]=8'b11111111;
memory[5677]=8'b11111111;
memory[5678]=8'b11111111;
memory[5679]=8'b11111111;
memory[5680]=8'b11111111;
memory[5681]=8'b11111111;
memory[5682]=8'b11111111;
memory[5683]=8'b11111111;
memory[5684]=8'b11111111;
memory[5685]=8'b11111111;
memory[5686]=8'b11111111;
memory[5687]=8'b11111111;
memory[5688]=8'b11111111;
memory[5689]=8'b11111111;
memory[5690]=8'b11111111;
memory[5691]=8'b11111111;
memory[5692]=8'b11100000;
memory[5693]=8'b11000011;
memory[5694]=8'b11111111;
memory[5695]=8'b11111111;
memory[5696]=8'b11111111;
memory[5697]=8'b11111111;
memory[5698]=8'b11111111;
memory[5699]=8'b11111111;
memory[5700]=8'b11111111;
memory[5701]=8'b11111111;
memory[5702]=8'b11111111;
memory[5703]=8'b11111111;
memory[5704]=8'b11111111;
memory[5705]=8'b11111111;
memory[5706]=8'b11111111;
memory[5707]=8'b11111100;
memory[5708]=8'b01110011;
memory[5709]=8'b11111111;
memory[5710]=8'b11111111;
memory[5711]=8'b11111111;
memory[5712]=8'b11111111;
memory[5713]=8'b11111111;
memory[5714]=8'b11111111;
memory[5715]=8'b11111111;
memory[5716]=8'b11111111;
memory[5717]=8'b11111111;
memory[5718]=8'b11111111;
memory[5719]=8'b11111111;
memory[5720]=8'b11111111;
memory[5721]=8'b11111111;
memory[5722]=8'b11111111;
memory[5723]=8'b11111111;
memory[5724]=8'b11111111;
memory[5725]=8'b11111111;
memory[5726]=8'b11111111;
memory[5727]=8'b11111111;
memory[5728]=8'b11111111;
memory[5729]=8'b11111111;
memory[5730]=8'b11111111;
memory[5731]=8'b11111111;
memory[5732]=8'b11110000;
memory[5733]=8'b11000011;
memory[5734]=8'b11111111;
memory[5735]=8'b11111111;
memory[5736]=8'b11111111;
memory[5737]=8'b11111111;
memory[5738]=8'b11111111;
memory[5739]=8'b11111111;
memory[5740]=8'b11111111;
memory[5741]=8'b11111111;
memory[5742]=8'b11111111;
memory[5743]=8'b11111111;
memory[5744]=8'b11111111;
memory[5745]=8'b11111111;
memory[5746]=8'b11111111;
memory[5747]=8'b11111100;
memory[5748]=8'b01110011;
memory[5749]=8'b11111111;
memory[5750]=8'b11111111;
memory[5751]=8'b11111111;
memory[5752]=8'b11111111;
memory[5753]=8'b11111111;
memory[5754]=8'b11111111;
memory[5755]=8'b11111111;
memory[5756]=8'b11111111;
memory[5757]=8'b11111111;
memory[5758]=8'b11111111;
memory[5759]=8'b11111111;
memory[5760]=8'b11111111;
memory[5761]=8'b11111111;
memory[5762]=8'b11111111;
memory[5763]=8'b11111111;
memory[5764]=8'b11111111;
memory[5765]=8'b11111111;
memory[5766]=8'b11111111;
memory[5767]=8'b11111111;
memory[5768]=8'b11111111;
memory[5769]=8'b11111111;
memory[5770]=8'b11111111;
memory[5771]=8'b11111111;
memory[5772]=8'b11110000;
memory[5773]=8'b11000011;
memory[5774]=8'b11111111;
memory[5775]=8'b11111111;
memory[5776]=8'b11111111;
memory[5777]=8'b11111111;
memory[5778]=8'b11111111;
memory[5779]=8'b11111111;
memory[5780]=8'b11111111;
memory[5781]=8'b11111111;
memory[5782]=8'b11111111;
memory[5783]=8'b11111111;
memory[5784]=8'b11111111;
memory[5785]=8'b11111111;
memory[5786]=8'b11111111;
memory[5787]=8'b11111100;
memory[5788]=8'b01110011;
memory[5789]=8'b11111111;
memory[5790]=8'b11111111;
memory[5791]=8'b11111111;
memory[5792]=8'b11111111;
memory[5793]=8'b11111111;
memory[5794]=8'b11111111;
memory[5795]=8'b11111111;
memory[5796]=8'b11111111;
memory[5797]=8'b11111111;
memory[5798]=8'b11111111;
memory[5799]=8'b11111111;
memory[5800]=8'b11111111;
memory[5801]=8'b11111111;
memory[5802]=8'b11111111;
memory[5803]=8'b11111111;
memory[5804]=8'b11111111;
memory[5805]=8'b11111111;
memory[5806]=8'b11111111;
memory[5807]=8'b11111111;
memory[5808]=8'b11111111;
memory[5809]=8'b11111111;
memory[5810]=8'b11111111;
memory[5811]=8'b11111111;
memory[5812]=8'b11111000;
memory[5813]=8'b01100011;
memory[5814]=8'b11111111;
memory[5815]=8'b11111111;
memory[5816]=8'b11111111;
memory[5817]=8'b11111111;
memory[5818]=8'b11111111;
memory[5819]=8'b11111111;
memory[5820]=8'b11111111;
memory[5821]=8'b11111111;
memory[5822]=8'b11111111;
memory[5823]=8'b11111111;
memory[5824]=8'b11111111;
memory[5825]=8'b11111111;
memory[5826]=8'b11111111;
memory[5827]=8'b11111110;
memory[5828]=8'b00111001;
memory[5829]=8'b11111111;
memory[5830]=8'b11111111;
memory[5831]=8'b11111111;
memory[5832]=8'b11111111;
memory[5833]=8'b11111111;
memory[5834]=8'b11111111;
memory[5835]=8'b11111111;
memory[5836]=8'b11111111;
memory[5837]=8'b11111111;
memory[5838]=8'b11111111;
memory[5839]=8'b11111111;
memory[5840]=8'b11111111;
memory[5841]=8'b11111111;
memory[5842]=8'b11111111;
memory[5843]=8'b11111111;
memory[5844]=8'b11111111;
memory[5845]=8'b11111111;
memory[5846]=8'b11111111;
memory[5847]=8'b11111111;
memory[5848]=8'b11111111;
memory[5849]=8'b11111111;
memory[5850]=8'b11111111;
memory[5851]=8'b11111111;
memory[5852]=8'b11111000;
memory[5853]=8'b01100011;
memory[5854]=8'b11111111;
memory[5855]=8'b11111111;
memory[5856]=8'b11111111;
memory[5857]=8'b11111111;
memory[5858]=8'b11111111;
memory[5859]=8'b11111111;
memory[5860]=8'b11111111;
memory[5861]=8'b11111111;
memory[5862]=8'b11111111;
memory[5863]=8'b11111111;
memory[5864]=8'b11111111;
memory[5865]=8'b11111111;
memory[5866]=8'b11111111;
memory[5867]=8'b11111110;
memory[5868]=8'b00111001;
memory[5869]=8'b11111111;
memory[5870]=8'b11111111;
memory[5871]=8'b11111111;
memory[5872]=8'b11111111;
memory[5873]=8'b11111111;
memory[5874]=8'b11111111;
memory[5875]=8'b11111111;
memory[5876]=8'b11111111;
memory[5877]=8'b11111111;
memory[5878]=8'b11111111;
memory[5879]=8'b11111111;
memory[5880]=8'b11111111;
memory[5881]=8'b11111111;
memory[5882]=8'b11111111;
memory[5883]=8'b11111111;
memory[5884]=8'b11111111;
memory[5885]=8'b11111111;
memory[5886]=8'b11111111;
memory[5887]=8'b11111111;
memory[5888]=8'b11111111;
memory[5889]=8'b11111111;
memory[5890]=8'b11111111;
memory[5891]=8'b11111111;
memory[5892]=8'b11111100;
memory[5893]=8'b01110011;
memory[5894]=8'b11111111;
memory[5895]=8'b11111111;
memory[5896]=8'b11111111;
memory[5897]=8'b11111111;
memory[5898]=8'b11111111;
memory[5899]=8'b11111111;
memory[5900]=8'b11111111;
memory[5901]=8'b11111111;
memory[5902]=8'b11111111;
memory[5903]=8'b11111111;
memory[5904]=8'b11111001;
memory[5905]=8'b11111111;
memory[5906]=8'b11111111;
memory[5907]=8'b11111110;
memory[5908]=8'b00111001;
memory[5909]=8'b11111111;
memory[5910]=8'b11111111;
memory[5911]=8'b11111111;
memory[5912]=8'b11111111;
memory[5913]=8'b11111111;
memory[5914]=8'b11111111;
memory[5915]=8'b11111111;
memory[5916]=8'b11111111;
memory[5917]=8'b11111111;
memory[5918]=8'b11111111;
memory[5919]=8'b11111111;
memory[5920]=8'b11111111;
memory[5921]=8'b11111111;
memory[5922]=8'b11111111;
memory[5923]=8'b11111111;
memory[5924]=8'b11111111;
memory[5925]=8'b11111111;
memory[5926]=8'b11111111;
memory[5927]=8'b11111111;
memory[5928]=8'b11111111;
memory[5929]=8'b11111111;
memory[5930]=8'b11111111;
memory[5931]=8'b11111111;
memory[5932]=8'b11111100;
memory[5933]=8'b00110011;
memory[5934]=8'b11111111;
memory[5935]=8'b11111111;
memory[5936]=8'b11111111;
memory[5937]=8'b11111111;
memory[5938]=8'b11111111;
memory[5939]=8'b11111111;
memory[5940]=8'b11111111;
memory[5941]=8'b11111111;
memory[5942]=8'b11111111;
memory[5943]=8'b11111111;
memory[5944]=8'b11110000;
memory[5945]=8'b00111111;
memory[5946]=8'b11111111;
memory[5947]=8'b11111110;
memory[5948]=8'b00111001;
memory[5949]=8'b11111111;
memory[5950]=8'b11111111;
memory[5951]=8'b11111111;
memory[5952]=8'b11111111;
memory[5953]=8'b11111111;
memory[5954]=8'b11111111;
memory[5955]=8'b11111111;
memory[5956]=8'b11111111;
memory[5957]=8'b11111111;
memory[5958]=8'b11111111;
memory[5959]=8'b11111111;
memory[5960]=8'b11111111;
memory[5961]=8'b11111111;
memory[5962]=8'b11111111;
memory[5963]=8'b11111111;
memory[5964]=8'b11111111;
memory[5965]=8'b11111111;
memory[5966]=8'b11111111;
memory[5967]=8'b11111111;
memory[5968]=8'b11111111;
memory[5969]=8'b11111111;
memory[5970]=8'b11111111;
memory[5971]=8'b11111111;
memory[5972]=8'b11111110;
memory[5973]=8'b00111111;
memory[5974]=8'b11111111;
memory[5975]=8'b11111111;
memory[5976]=8'b11111111;
memory[5977]=8'b11111111;
memory[5978]=8'b11111111;
memory[5979]=8'b11111111;
memory[5980]=8'b11111111;
memory[5981]=8'b11111111;
memory[5982]=8'b11111111;
memory[5983]=8'b11111111;
memory[5984]=8'b11100001;
memory[5985]=8'b11111111;
memory[5986]=8'b11111111;
memory[5987]=8'b11111110;
memory[5988]=8'b00111000;
memory[5989]=8'b11111111;
memory[5990]=8'b11111111;
memory[5991]=8'b11111111;
memory[5992]=8'b11111111;
memory[5993]=8'b11111111;
memory[5994]=8'b11111111;
memory[5995]=8'b11111111;
memory[5996]=8'b11111111;
memory[5997]=8'b11111111;
memory[5998]=8'b11111111;
memory[5999]=8'b11111111;
memory[6000]=8'b11111111;
memory[6001]=8'b11111111;
memory[6002]=8'b11111111;
memory[6003]=8'b11111111;
memory[6004]=8'b11111111;
memory[6005]=8'b11111111;
memory[6006]=8'b11111111;
memory[6007]=8'b11111111;
memory[6008]=8'b11111111;
memory[6009]=8'b11111111;
memory[6010]=8'b11111111;
memory[6011]=8'b11111111;
memory[6012]=8'b11111110;
memory[6013]=8'b00011111;
memory[6014]=8'b11111111;
memory[6015]=8'b11111111;
memory[6016]=8'b11111111;
memory[6017]=8'b11111111;
memory[6018]=8'b11111111;
memory[6019]=8'b11111111;
memory[6020]=8'b11111111;
memory[6021]=8'b11111111;
memory[6022]=8'b11111111;
memory[6023]=8'b11111111;
memory[6024]=8'b11100111;
memory[6025]=8'b11111111;
memory[6026]=8'b11111111;
memory[6027]=8'b11111110;
memory[6028]=8'b00111000;
memory[6029]=8'b11111111;
memory[6030]=8'b11111111;
memory[6031]=8'b11111111;
memory[6032]=8'b11111111;
memory[6033]=8'b11111111;
memory[6034]=8'b11111111;
memory[6035]=8'b11111111;
memory[6036]=8'b11111111;
memory[6037]=8'b11111111;
memory[6038]=8'b11111111;
memory[6039]=8'b11111111;
memory[6040]=8'b11111111;
memory[6041]=8'b11111111;
memory[6042]=8'b11111111;
memory[6043]=8'b11111111;
memory[6044]=8'b11111111;
memory[6045]=8'b11111111;
memory[6046]=8'b11111111;
memory[6047]=8'b11111111;
memory[6048]=8'b11111111;
memory[6049]=8'b11111111;
memory[6050]=8'b11111111;
memory[6051]=8'b11111111;
memory[6052]=8'b11111111;
memory[6053]=8'b00001111;
memory[6054]=8'b11111111;
memory[6055]=8'b11111111;
memory[6056]=8'b11111111;
memory[6057]=8'b11111111;
memory[6058]=8'b11111111;
memory[6059]=8'b11111111;
memory[6060]=8'b11111111;
memory[6061]=8'b11111111;
memory[6062]=8'b11111111;
memory[6063]=8'b11111111;
memory[6064]=8'b11001111;
memory[6065]=8'b11111111;
memory[6066]=8'b11111111;
memory[6067]=8'b11111100;
memory[6068]=8'b00110000;
memory[6069]=8'b11111111;
memory[6070]=8'b11111111;
memory[6071]=8'b11111111;
memory[6072]=8'b11111111;
memory[6073]=8'b11111111;
memory[6074]=8'b11111111;
memory[6075]=8'b11111111;
memory[6076]=8'b11111111;
memory[6077]=8'b11111111;
memory[6078]=8'b11111111;
memory[6079]=8'b11111111;
memory[6080]=8'b11111111;
memory[6081]=8'b11111111;
memory[6082]=8'b11111111;
memory[6083]=8'b11111111;
memory[6084]=8'b11111111;
memory[6085]=8'b11111111;
memory[6086]=8'b11111111;
memory[6087]=8'b11111111;
memory[6088]=8'b11111111;
memory[6089]=8'b11111111;
memory[6090]=8'b11111111;
memory[6091]=8'b11111111;
memory[6092]=8'b11111111;
memory[6093]=8'b00001111;
memory[6094]=8'b11111111;
memory[6095]=8'b11111111;
memory[6096]=8'b11111111;
memory[6097]=8'b11111111;
memory[6098]=8'b11111111;
memory[6099]=8'b11111111;
memory[6100]=8'b11111111;
memory[6101]=8'b11111111;
memory[6102]=8'b11000011;
memory[6103]=8'b11111111;
memory[6104]=8'b11011111;
memory[6105]=8'b11111111;
memory[6106]=8'b11111111;
memory[6107]=8'b11111100;
memory[6108]=8'b00110000;
memory[6109]=8'b01111111;
memory[6110]=8'b11111111;
memory[6111]=8'b11111111;
memory[6112]=8'b11111111;
memory[6113]=8'b11111111;
memory[6114]=8'b11111111;
memory[6115]=8'b11111111;
memory[6116]=8'b11111111;
memory[6117]=8'b11111111;
memory[6118]=8'b11111111;
memory[6119]=8'b11111111;
memory[6120]=8'b11111111;
memory[6121]=8'b11111111;
memory[6122]=8'b11111111;
memory[6123]=8'b11111111;
memory[6124]=8'b11111111;
memory[6125]=8'b11111111;
memory[6126]=8'b11111111;
memory[6127]=8'b11111111;
memory[6128]=8'b11111111;
memory[6129]=8'b11111111;
memory[6130]=8'b11111111;
memory[6131]=8'b11111111;
memory[6132]=8'b11111111;
memory[6133]=8'b10001111;
memory[6134]=8'b11111111;
memory[6135]=8'b11111111;
memory[6136]=8'b11111111;
memory[6137]=8'b11111111;
memory[6138]=8'b11111111;
memory[6139]=8'b11111111;
memory[6140]=8'b11111111;
memory[6141]=8'b11111111;
memory[6142]=8'b11111111;
memory[6143]=8'b11111111;
memory[6144]=8'b11111111;
memory[6145]=8'b11111111;
memory[6146]=8'b11111111;
memory[6147]=8'b11111100;
memory[6148]=8'b00110000;
memory[6149]=8'b11111111;
memory[6150]=8'b11111111;
memory[6151]=8'b11111111;
memory[6152]=8'b11111111;
memory[6153]=8'b11111111;
memory[6154]=8'b11111111;
memory[6155]=8'b11111111;
memory[6156]=8'b11111111;
memory[6157]=8'b11111111;
memory[6158]=8'b11111111;
memory[6159]=8'b11111111;
memory[6160]=8'b11111111;
memory[6161]=8'b11111111;
memory[6162]=8'b11111111;
memory[6163]=8'b11111111;
memory[6164]=8'b11111111;
memory[6165]=8'b11111111;
memory[6166]=8'b11111111;
memory[6167]=8'b11111111;
memory[6168]=8'b11111111;
memory[6169]=8'b11111111;
memory[6170]=8'b11111111;
memory[6171]=8'b11111111;
memory[6172]=8'b11111111;
memory[6173]=8'b10000111;
memory[6174]=8'b11111111;
memory[6175]=8'b11111111;
memory[6176]=8'b11111111;
memory[6177]=8'b11111111;
memory[6178]=8'b11111111;
memory[6179]=8'b11111111;
memory[6180]=8'b11111111;
memory[6181]=8'b11111111;
memory[6182]=8'b11111111;
memory[6183]=8'b11111111;
memory[6184]=8'b11111111;
memory[6185]=8'b11111111;
memory[6186]=8'b11111111;
memory[6187]=8'b11111100;
memory[6188]=8'b00100000;
memory[6189]=8'b11111111;
memory[6190]=8'b11111111;
memory[6191]=8'b11111111;
memory[6192]=8'b11111111;
memory[6193]=8'b11111111;
memory[6194]=8'b11111111;
memory[6195]=8'b11111111;
memory[6196]=8'b11111111;
memory[6197]=8'b11111111;
memory[6198]=8'b11111111;
memory[6199]=8'b11111111;
memory[6200]=8'b11111111;
memory[6201]=8'b11111111;
memory[6202]=8'b11111111;
memory[6203]=8'b11111111;
memory[6204]=8'b11111111;
memory[6205]=8'b11111111;
memory[6206]=8'b11111111;
memory[6207]=8'b11111111;
memory[6208]=8'b11111111;
memory[6209]=8'b11111111;
memory[6210]=8'b11111111;
memory[6211]=8'b11111111;
memory[6212]=8'b11111111;
memory[6213]=8'b11000111;
memory[6214]=8'b11111111;
memory[6215]=8'b11111111;
memory[6216]=8'b11111111;
memory[6217]=8'b11111111;
memory[6218]=8'b11111111;
memory[6219]=8'b11111111;
memory[6220]=8'b11111111;
memory[6221]=8'b11111111;
memory[6222]=8'b11111110;
memory[6223]=8'b11111111;
memory[6224]=8'b11111111;
memory[6225]=8'b11111111;
memory[6226]=8'b11111111;
memory[6227]=8'b11111110;
memory[6228]=8'b00100001;
memory[6229]=8'b11111111;
memory[6230]=8'b11111111;
memory[6231]=8'b11111111;
memory[6232]=8'b11111111;
memory[6233]=8'b11111111;
memory[6234]=8'b11111111;
memory[6235]=8'b11111111;
memory[6236]=8'b11111111;
memory[6237]=8'b11111111;
memory[6238]=8'b11111111;
memory[6239]=8'b11111111;
memory[6240]=8'b11111111;
memory[6241]=8'b11111111;
memory[6242]=8'b11111111;
memory[6243]=8'b11111111;
memory[6244]=8'b11111111;
memory[6245]=8'b11111111;
memory[6246]=8'b11111111;
memory[6247]=8'b11111111;
memory[6248]=8'b11111111;
memory[6249]=8'b11111111;
memory[6250]=8'b11111111;
memory[6251]=8'b11111111;
memory[6252]=8'b11111111;
memory[6253]=8'b11000111;
memory[6254]=8'b11111111;
memory[6255]=8'b11111111;
memory[6256]=8'b11111111;
memory[6257]=8'b11111111;
memory[6258]=8'b11111111;
memory[6259]=8'b11111111;
memory[6260]=8'b11111111;
memory[6261]=8'b11111111;
memory[6262]=8'b11111100;
memory[6263]=8'b00011111;
memory[6264]=8'b11111100;
memory[6265]=8'b11111111;
memory[6266]=8'b11111111;
memory[6267]=8'b11111110;
memory[6268]=8'b01000011;
memory[6269]=8'b11111111;
memory[6270]=8'b11111111;
memory[6271]=8'b11111111;
memory[6272]=8'b11111111;
memory[6273]=8'b11111111;
memory[6274]=8'b11111111;
memory[6275]=8'b11111111;
memory[6276]=8'b11111111;
memory[6277]=8'b11111111;
memory[6278]=8'b11111111;
memory[6279]=8'b11111111;
memory[6280]=8'b11111111;
memory[6281]=8'b11111111;
memory[6282]=8'b11111111;
memory[6283]=8'b11111111;
memory[6284]=8'b11111111;
memory[6285]=8'b11111111;
memory[6286]=8'b11111111;
memory[6287]=8'b11111111;
memory[6288]=8'b11111111;
memory[6289]=8'b11111111;
memory[6290]=8'b11111111;
memory[6291]=8'b11111111;
memory[6292]=8'b11111111;
memory[6293]=8'b11100011;
memory[6294]=8'b11111111;
memory[6295]=8'b11111111;
memory[6296]=8'b11111111;
memory[6297]=8'b11111111;
memory[6298]=8'b11111111;
memory[6299]=8'b11111111;
memory[6300]=8'b11111111;
memory[6301]=8'b11111111;
memory[6302]=8'b11111111;
memory[6303]=8'b00000111;
memory[6304]=8'b11111101;
memory[6305]=8'b11111111;
memory[6306]=8'b11111111;
memory[6307]=8'b11111110;
memory[6308]=8'b01000011;
memory[6309]=8'b11111111;
memory[6310]=8'b11111111;
memory[6311]=8'b11111111;
memory[6312]=8'b11111111;
memory[6313]=8'b11111111;
memory[6314]=8'b11111111;
memory[6315]=8'b11111111;
memory[6316]=8'b11111111;
memory[6317]=8'b11111111;
memory[6318]=8'b11111111;
memory[6319]=8'b11111111;
memory[6320]=8'b11111111;
memory[6321]=8'b11111111;
memory[6322]=8'b11111111;
memory[6323]=8'b11111111;
memory[6324]=8'b11111111;
memory[6325]=8'b11111111;
memory[6326]=8'b11111111;
memory[6327]=8'b11111111;
memory[6328]=8'b11111111;
memory[6329]=8'b11111111;
memory[6330]=8'b11111111;
memory[6331]=8'b11111111;
memory[6332]=8'b11111111;
memory[6333]=8'b11100011;
memory[6334]=8'b11111111;
memory[6335]=8'b11111111;
memory[6336]=8'b11111111;
memory[6337]=8'b11111111;
memory[6338]=8'b11111111;
memory[6339]=8'b11111111;
memory[6340]=8'b11111111;
memory[6341]=8'b11111111;
memory[6342]=8'b11111111;
memory[6343]=8'b11000011;
memory[6344]=8'b11111111;
memory[6345]=8'b11111111;
memory[6346]=8'b11111111;
memory[6347]=8'b11111110;
memory[6348]=8'b01000111;
memory[6349]=8'b11111111;
memory[6350]=8'b11111111;
memory[6351]=8'b11111111;
memory[6352]=8'b11111111;
memory[6353]=8'b11111111;
memory[6354]=8'b11111111;
memory[6355]=8'b11111111;
memory[6356]=8'b11111111;
memory[6357]=8'b11111111;
memory[6358]=8'b11111111;
memory[6359]=8'b11111111;
memory[6360]=8'b11111111;
memory[6361]=8'b11111111;
memory[6362]=8'b11111111;
memory[6363]=8'b11111111;
memory[6364]=8'b11111111;
memory[6365]=8'b11111111;
memory[6366]=8'b11111111;
memory[6367]=8'b11111111;
memory[6368]=8'b11111111;
memory[6369]=8'b11111111;
memory[6370]=8'b11111111;
memory[6371]=8'b11111111;
memory[6372]=8'b11111111;
memory[6373]=8'b11100011;
memory[6374]=8'b11111111;
memory[6375]=8'b11111111;
memory[6376]=8'b11111111;
memory[6377]=8'b11111111;
memory[6378]=8'b11111111;
memory[6379]=8'b11111111;
memory[6380]=8'b11111111;
memory[6381]=8'b11111111;
memory[6382]=8'b11111111;
memory[6383]=8'b00000000;
memory[6384]=8'b11111111;
memory[6385]=8'b11111111;
memory[6386]=8'b11111111;
memory[6387]=8'b11111100;
memory[6388]=8'b00000111;
memory[6389]=8'b11111111;
memory[6390]=8'b11111111;
memory[6391]=8'b11111111;
memory[6392]=8'b11111111;
memory[6393]=8'b11111111;
memory[6394]=8'b11111111;
memory[6395]=8'b11111111;
memory[6396]=8'b11111111;
memory[6397]=8'b11111111;
memory[6398]=8'b11111111;
memory[6399]=8'b11111111;
memory[6400]=8'b11111111;
memory[6401]=8'b11111111;
memory[6402]=8'b11111111;
memory[6403]=8'b11111111;
memory[6404]=8'b11111111;
memory[6405]=8'b11111111;
memory[6406]=8'b11111111;
memory[6407]=8'b11111111;
memory[6408]=8'b11111111;
memory[6409]=8'b11111111;
memory[6410]=8'b11111111;
memory[6411]=8'b11111111;
memory[6412]=8'b11111111;
memory[6413]=8'b11110001;
memory[6414]=8'b11111111;
memory[6415]=8'b11111111;
memory[6416]=8'b11111111;
memory[6417]=8'b11111111;
memory[6418]=8'b11111111;
memory[6419]=8'b11111111;
memory[6420]=8'b11111111;
memory[6421]=8'b11111111;
memory[6422]=8'b11111111;
memory[6423]=8'b11000000;
memory[6424]=8'b01111111;
memory[6425]=8'b11111111;
memory[6426]=8'b11111111;
memory[6427]=8'b11111111;
memory[6428]=8'b10001111;
memory[6429]=8'b11111111;
memory[6430]=8'b11111111;
memory[6431]=8'b11111111;
memory[6432]=8'b11111111;
memory[6433]=8'b11111111;
memory[6434]=8'b11111111;
memory[6435]=8'b11111111;
memory[6436]=8'b11111111;
memory[6437]=8'b11111111;
memory[6438]=8'b11111111;
memory[6439]=8'b11111111;
memory[6440]=8'b11111111;
memory[6441]=8'b11111111;
memory[6442]=8'b11111111;
memory[6443]=8'b11111111;
memory[6444]=8'b11111111;
memory[6445]=8'b11111111;
memory[6446]=8'b11111111;
memory[6447]=8'b11111111;
memory[6448]=8'b11111111;
memory[6449]=8'b11111111;
memory[6450]=8'b11111111;
memory[6451]=8'b11111111;
memory[6452]=8'b11111111;
memory[6453]=8'b11110001;
memory[6454]=8'b11111111;
memory[6455]=8'b11111111;
memory[6456]=8'b11111111;
memory[6457]=8'b11111111;
memory[6458]=8'b11111111;
memory[6459]=8'b11111111;
memory[6460]=8'b11111111;
memory[6461]=8'b11111111;
memory[6462]=8'b11111111;
memory[6463]=8'b11111100;
memory[6464]=8'b01111111;
memory[6465]=8'b11111111;
memory[6466]=8'b11111111;
memory[6467]=8'b11111111;
memory[6468]=8'b10001111;
memory[6469]=8'b11111111;
memory[6470]=8'b11111111;
memory[6471]=8'b11111111;
memory[6472]=8'b11111111;
memory[6473]=8'b11111111;
memory[6474]=8'b11111111;
memory[6475]=8'b11111111;
memory[6476]=8'b11111111;
memory[6477]=8'b11111111;
memory[6478]=8'b11111111;
memory[6479]=8'b11111111;
memory[6480]=8'b11111111;
memory[6481]=8'b11111111;
memory[6482]=8'b11111111;
memory[6483]=8'b11111111;
memory[6484]=8'b11111111;
memory[6485]=8'b11111111;
memory[6486]=8'b11111111;
memory[6487]=8'b11111111;
memory[6488]=8'b11111111;
memory[6489]=8'b11111111;
memory[6490]=8'b11111111;
memory[6491]=8'b11111111;
memory[6492]=8'b11111111;
memory[6493]=8'b11111001;
memory[6494]=8'b11111111;
memory[6495]=8'b11111111;
memory[6496]=8'b11111111;
memory[6497]=8'b11111111;
memory[6498]=8'b11111111;
memory[6499]=8'b11111111;
memory[6500]=8'b11111111;
memory[6501]=8'b11111111;
memory[6502]=8'b11111111;
memory[6503]=8'b11111111;
memory[6504]=8'b00111111;
memory[6505]=8'b11111111;
memory[6506]=8'b11111111;
memory[6507]=8'b11111111;
memory[6508]=8'b00011111;
memory[6509]=8'b11111111;
memory[6510]=8'b11111111;
memory[6511]=8'b11111111;
memory[6512]=8'b11111111;
memory[6513]=8'b11111111;
memory[6514]=8'b11111111;
memory[6515]=8'b11111111;
memory[6516]=8'b11111111;
memory[6517]=8'b11111111;
memory[6518]=8'b11111111;
memory[6519]=8'b11111111;
memory[6520]=8'b11111111;
memory[6521]=8'b11111111;
memory[6522]=8'b11111111;
memory[6523]=8'b11111111;
memory[6524]=8'b11111111;
memory[6525]=8'b11111111;
memory[6526]=8'b11111111;
memory[6527]=8'b11111111;
memory[6528]=8'b11111111;
memory[6529]=8'b11111111;
memory[6530]=8'b11111111;
memory[6531]=8'b11111111;
memory[6532]=8'b11111111;
memory[6533]=8'b11111001;
memory[6534]=8'b11111111;
memory[6535]=8'b11111111;
memory[6536]=8'b11111111;
memory[6537]=8'b11111111;
memory[6538]=8'b11111111;
memory[6539]=8'b11111111;
memory[6540]=8'b11111111;
memory[6541]=8'b11111111;
memory[6542]=8'b11111111;
memory[6543]=8'b11111111;
memory[6544]=8'b10011111;
memory[6545]=8'b11111111;
memory[6546]=8'b11111111;
memory[6547]=8'b11111111;
memory[6548]=8'b00011111;
memory[6549]=8'b11111111;
memory[6550]=8'b11111111;
memory[6551]=8'b11111111;
memory[6552]=8'b11111111;
memory[6553]=8'b11111111;
memory[6554]=8'b11111111;
memory[6555]=8'b11111111;
memory[6556]=8'b11111111;
memory[6557]=8'b11111111;
memory[6558]=8'b11111111;
memory[6559]=8'b11111111;
memory[6560]=8'b11111111;
memory[6561]=8'b11111111;
memory[6562]=8'b11111111;
memory[6563]=8'b11111111;
memory[6564]=8'b11111111;
memory[6565]=8'b11111111;
memory[6566]=8'b11111111;
memory[6567]=8'b11111111;
memory[6568]=8'b11111111;
memory[6569]=8'b11111111;
memory[6570]=8'b11111111;
memory[6571]=8'b11111111;
memory[6572]=8'b11111111;
memory[6573]=8'b11111000;
memory[6574]=8'b11111111;
memory[6575]=8'b11111111;
memory[6576]=8'b11111111;
memory[6577]=8'b11111111;
memory[6578]=8'b11111111;
memory[6579]=8'b11111111;
memory[6580]=8'b11111111;
memory[6581]=8'b11111111;
memory[6582]=8'b11111111;
memory[6583]=8'b11111111;
memory[6584]=8'b10011111;
memory[6585]=8'b11111111;
memory[6586]=8'b11111111;
memory[6587]=8'b11111111;
memory[6588]=8'b00111111;
memory[6589]=8'b11111111;
memory[6590]=8'b11111111;
memory[6591]=8'b11111111;
memory[6592]=8'b11111111;
memory[6593]=8'b11111111;
memory[6594]=8'b11111111;
memory[6595]=8'b11111111;
memory[6596]=8'b11111111;
memory[6597]=8'b11111111;
memory[6598]=8'b11111111;
memory[6599]=8'b11111111;
memory[6600]=8'b11111111;
memory[6601]=8'b11111111;
memory[6602]=8'b11111111;
memory[6603]=8'b11111111;
memory[6604]=8'b11111111;
memory[6605]=8'b11111111;
memory[6606]=8'b11111111;
memory[6607]=8'b11111111;
memory[6608]=8'b11111111;
memory[6609]=8'b11111111;
memory[6610]=8'b11111111;
memory[6611]=8'b11111111;
memory[6612]=8'b11111111;
memory[6613]=8'b11111100;
memory[6614]=8'b11111111;
memory[6615]=8'b11111111;
memory[6616]=8'b11111111;
memory[6617]=8'b11111111;
memory[6618]=8'b11111111;
memory[6619]=8'b11111111;
memory[6620]=8'b11111111;
memory[6621]=8'b11111111;
memory[6622]=8'b11111111;
memory[6623]=8'b11111111;
memory[6624]=8'b10011111;
memory[6625]=8'b11111111;
memory[6626]=8'b11111111;
memory[6627]=8'b11111110;
memory[6628]=8'b00111111;
memory[6629]=8'b11111111;
memory[6630]=8'b11111111;
memory[6631]=8'b11111111;
memory[6632]=8'b11111111;
memory[6633]=8'b11111111;
memory[6634]=8'b11111111;
memory[6635]=8'b11111111;
memory[6636]=8'b11111111;
memory[6637]=8'b11111111;
memory[6638]=8'b11111111;
memory[6639]=8'b11111111;
memory[6640]=8'b11111111;
memory[6641]=8'b11111111;
memory[6642]=8'b11111111;
memory[6643]=8'b11111111;
memory[6644]=8'b11111111;
memory[6645]=8'b11111111;
memory[6646]=8'b11111111;
memory[6647]=8'b11111111;
memory[6648]=8'b11111111;
memory[6649]=8'b11111111;
memory[6650]=8'b11111111;
memory[6651]=8'b11111111;
memory[6652]=8'b11111111;
memory[6653]=8'b11111100;
memory[6654]=8'b11111111;
memory[6655]=8'b11111111;
memory[6656]=8'b11111111;
memory[6657]=8'b11111111;
memory[6658]=8'b11111111;
memory[6659]=8'b11111111;
memory[6660]=8'b11111111;
memory[6661]=8'b11111111;
memory[6662]=8'b11111111;
memory[6663]=8'b11111111;
memory[6664]=8'b00111111;
memory[6665]=8'b11110000;
memory[6666]=8'b00000111;
memory[6667]=8'b11111110;
memory[6668]=8'b01111111;
memory[6669]=8'b11111111;
memory[6670]=8'b11111111;
memory[6671]=8'b11111111;
memory[6672]=8'b11111111;
memory[6673]=8'b11111111;
memory[6674]=8'b11111111;
memory[6675]=8'b11111111;
memory[6676]=8'b11111111;
memory[6677]=8'b11111111;
memory[6678]=8'b11111111;
memory[6679]=8'b11111111;
memory[6680]=8'b11111111;
memory[6681]=8'b11111111;
memory[6682]=8'b11111111;
memory[6683]=8'b11111111;
memory[6684]=8'b11111111;
memory[6685]=8'b11111111;
memory[6686]=8'b11111111;
memory[6687]=8'b11111111;
memory[6688]=8'b11111111;
memory[6689]=8'b11111111;
memory[6690]=8'b11111111;
memory[6691]=8'b11111111;
memory[6692]=8'b11111111;
memory[6693]=8'b11111100;
memory[6694]=8'b11111111;
memory[6695]=8'b11111111;
memory[6696]=8'b11111111;
memory[6697]=8'b11111111;
memory[6698]=8'b11111111;
memory[6699]=8'b11111111;
memory[6700]=8'b11111000;
memory[6701]=8'b11111111;
memory[6702]=8'b11111111;
memory[6703]=8'b11111000;
memory[6704]=8'b01111111;
memory[6705]=8'b10000111;
memory[6706]=8'b11111111;
memory[6707]=8'b11111110;
memory[6708]=8'b01111111;
memory[6709]=8'b11111111;
memory[6710]=8'b11111111;
memory[6711]=8'b11111111;
memory[6712]=8'b11111111;
memory[6713]=8'b11111111;
memory[6714]=8'b11111111;
memory[6715]=8'b11111111;
memory[6716]=8'b11111111;
memory[6717]=8'b11111111;
memory[6718]=8'b11111111;
memory[6719]=8'b11111111;
memory[6720]=8'b11111111;
memory[6721]=8'b11111111;
memory[6722]=8'b11111111;
memory[6723]=8'b11111111;
memory[6724]=8'b11111111;
memory[6725]=8'b11111111;
memory[6726]=8'b11111111;
memory[6727]=8'b11111111;
memory[6728]=8'b11111111;
memory[6729]=8'b11111111;
memory[6730]=8'b11111111;
memory[6731]=8'b11111111;
memory[6732]=8'b11111111;
memory[6733]=8'b11101110;
memory[6734]=8'b01111111;
memory[6735]=8'b11111111;
memory[6736]=8'b11111111;
memory[6737]=8'b11111111;
memory[6738]=8'b11111111;
memory[6739]=8'b11111111;
memory[6740]=8'b11111111;
memory[6741]=8'b10000000;
memory[6742]=8'b00001110;
memory[6743]=8'b00000011;
memory[6744]=8'b11111100;
memory[6745]=8'b01111111;
memory[6746]=8'b11111111;
memory[6747]=8'b11111100;
memory[6748]=8'b11111111;
memory[6749]=8'b11111111;
memory[6750]=8'b11111111;
memory[6751]=8'b11111111;
memory[6752]=8'b11111111;
memory[6753]=8'b11111111;
memory[6754]=8'b11111111;
memory[6755]=8'b11111111;
memory[6756]=8'b11111111;
memory[6757]=8'b11111111;
memory[6758]=8'b11111111;
memory[6759]=8'b11111111;
memory[6760]=8'b11111111;
memory[6761]=8'b11111111;
memory[6762]=8'b11111111;
memory[6763]=8'b11111111;
memory[6764]=8'b11111111;
memory[6765]=8'b11111111;
memory[6766]=8'b11111111;
memory[6767]=8'b11111111;
memory[6768]=8'b11111111;
memory[6769]=8'b11111111;
memory[6770]=8'b11111111;
memory[6771]=8'b11111111;
memory[6772]=8'b11111111;
memory[6773]=8'b11100110;
memory[6774]=8'b01111111;
memory[6775]=8'b11111111;
memory[6776]=8'b11111111;
memory[6777]=8'b11111111;
memory[6778]=8'b11111111;
memory[6779]=8'b11111111;
memory[6780]=8'b11111111;
memory[6781]=8'b11111111;
memory[6782]=8'b11000001;
memory[6783]=8'b11111111;
memory[6784]=8'b11000111;
memory[6785]=8'b11111111;
memory[6786]=8'b11111111;
memory[6787]=8'b11111100;
memory[6788]=8'b11111111;
memory[6789]=8'b11111111;
memory[6790]=8'b11111111;
memory[6791]=8'b11111111;
memory[6792]=8'b11111111;
memory[6793]=8'b11111111;
memory[6794]=8'b11111111;
memory[6795]=8'b11111111;
memory[6796]=8'b11111111;
memory[6797]=8'b11111111;
memory[6798]=8'b11111111;
memory[6799]=8'b11111111;
memory[6800]=8'b11111111;
memory[6801]=8'b11111111;
memory[6802]=8'b11111111;
memory[6803]=8'b11111111;
memory[6804]=8'b11111111;
memory[6805]=8'b11111111;
memory[6806]=8'b11111111;
memory[6807]=8'b11111111;
memory[6808]=8'b11111111;
memory[6809]=8'b11111111;
memory[6810]=8'b11111111;
memory[6811]=8'b11111111;
memory[6812]=8'b11111111;
memory[6813]=8'b11100110;
memory[6814]=8'b01111111;
memory[6815]=8'b11111111;
memory[6816]=8'b11111111;
memory[6817]=8'b11111111;
memory[6818]=8'b11111111;
memory[6819]=8'b11111111;
memory[6820]=8'b11111111;
memory[6821]=8'b11111111;
memory[6822]=8'b11111111;
memory[6823]=8'b11111100;
memory[6824]=8'b01111111;
memory[6825]=8'b11111111;
memory[6826]=8'b11111111;
memory[6827]=8'b11111101;
memory[6828]=8'b11111111;
memory[6829]=8'b11111111;
memory[6830]=8'b11111111;
memory[6831]=8'b11111111;
memory[6832]=8'b11111111;
memory[6833]=8'b11111111;
memory[6834]=8'b11111111;
memory[6835]=8'b11111111;
memory[6836]=8'b11111111;
memory[6837]=8'b11111111;
memory[6838]=8'b11111111;
memory[6839]=8'b11111111;
memory[6840]=8'b11111111;
memory[6841]=8'b11111111;
memory[6842]=8'b11111111;
memory[6843]=8'b11111111;
memory[6844]=8'b11111111;
memory[6845]=8'b11111111;
memory[6846]=8'b11111111;
memory[6847]=8'b11111111;
memory[6848]=8'b11111111;
memory[6849]=8'b11111111;
memory[6850]=8'b11111111;
memory[6851]=8'b11111111;
memory[6852]=8'b11111111;
memory[6853]=8'b11110110;
memory[6854]=8'b00111111;
memory[6855]=8'b11111111;
memory[6856]=8'b11111111;
memory[6857]=8'b11111111;
memory[6858]=8'b11111111;
memory[6859]=8'b11111111;
memory[6860]=8'b11111111;
memory[6861]=8'b11111111;
memory[6862]=8'b11111111;
memory[6863]=8'b11111111;
memory[6864]=8'b11111111;
memory[6865]=8'b11111111;
memory[6866]=8'b11111111;
memory[6867]=8'b11111101;
memory[6868]=8'b11111111;
memory[6869]=8'b11111100;
memory[6870]=8'b11111111;
memory[6871]=8'b11111111;
memory[6872]=8'b11111111;
memory[6873]=8'b11111111;
memory[6874]=8'b11111111;
memory[6875]=8'b11111111;
memory[6876]=8'b11111111;
memory[6877]=8'b11111111;
memory[6878]=8'b11111111;
memory[6879]=8'b11111111;
memory[6880]=8'b11111111;
memory[6881]=8'b11111111;
memory[6882]=8'b11111111;
memory[6883]=8'b11111111;
memory[6884]=8'b11111111;
memory[6885]=8'b11111111;
memory[6886]=8'b11111111;
memory[6887]=8'b11111111;
memory[6888]=8'b11111111;
memory[6889]=8'b11111111;
memory[6890]=8'b11111111;
memory[6891]=8'b11111111;
memory[6892]=8'b11111111;
memory[6893]=8'b11100110;
memory[6894]=8'b00111111;
memory[6895]=8'b11111111;
memory[6896]=8'b11111111;
memory[6897]=8'b10000000;
memory[6898]=8'b00000011;
memory[6899]=8'b11111111;
memory[6900]=8'b11111111;
memory[6901]=8'b11111111;
memory[6902]=8'b11111111;
memory[6903]=8'b11111111;
memory[6904]=8'b11111111;
memory[6905]=8'b11111111;
memory[6906]=8'b11111111;
memory[6907]=8'b11111001;
memory[6908]=8'b11111111;
memory[6909]=8'b11100000;
memory[6910]=8'b00001111;
memory[6911]=8'b11111111;
memory[6912]=8'b11111111;
memory[6913]=8'b11111111;
memory[6914]=8'b11111111;
memory[6915]=8'b11111111;
memory[6916]=8'b11111111;
memory[6917]=8'b11111111;
memory[6918]=8'b11111111;
memory[6919]=8'b11111111;
memory[6920]=8'b11111111;
memory[6921]=8'b11111111;
memory[6922]=8'b11111111;
memory[6923]=8'b11111111;
memory[6924]=8'b11111111;
memory[6925]=8'b11111111;
memory[6926]=8'b11111111;
memory[6927]=8'b11111111;
memory[6928]=8'b11111111;
memory[6929]=8'b11111111;
memory[6930]=8'b11111111;
memory[6931]=8'b11111111;
memory[6932]=8'b11111111;
memory[6933]=8'b11100011;
memory[6934]=8'b00111111;
memory[6935]=8'b11111111;
memory[6936]=8'b11111111;
memory[6937]=8'b11111111;
memory[6938]=8'b00000000;
memory[6939]=8'b00000011;
memory[6940]=8'b11111111;
memory[6941]=8'b11111111;
memory[6942]=8'b11111111;
memory[6943]=8'b11111111;
memory[6944]=8'b11111111;
memory[6945]=8'b11111111;
memory[6946]=8'b11111111;
memory[6947]=8'b11111000;
memory[6948]=8'b11111111;
memory[6949]=8'b11111111;
memory[6950]=8'b10000001;
memory[6951]=8'b11111111;
memory[6952]=8'b11111111;
memory[6953]=8'b11111111;
memory[6954]=8'b11111111;
memory[6955]=8'b11111111;
memory[6956]=8'b11111111;
memory[6957]=8'b11111111;
memory[6958]=8'b11111111;
memory[6959]=8'b11111111;
memory[6960]=8'b11111111;
memory[6961]=8'b11111111;
memory[6962]=8'b11111111;
memory[6963]=8'b11111111;
memory[6964]=8'b11111111;
memory[6965]=8'b11111111;
memory[6966]=8'b11111111;
memory[6967]=8'b11111100;
memory[6968]=8'b00000000;
memory[6969]=8'b01111111;
memory[6970]=8'b11111111;
memory[6971]=8'b11111111;
memory[6972]=8'b11111111;
memory[6973]=8'b11110001;
memory[6974]=8'b00011111;
memory[6975]=8'b11111111;
memory[6976]=8'b11111111;
memory[6977]=8'b11111111;
memory[6978]=8'b11111100;
memory[6979]=8'b00000000;
memory[6980]=8'b00111111;
memory[6981]=8'b11111111;
memory[6982]=8'b11111111;
memory[6983]=8'b11111111;
memory[6984]=8'b10001111;
memory[6985]=8'b11111111;
memory[6986]=8'b11111111;
memory[6987]=8'b11111000;
memory[6988]=8'b11111111;
memory[6989]=8'b11111111;
memory[6990]=8'b11111000;
memory[6991]=8'b00000000;
memory[6992]=8'b01111111;
memory[6993]=8'b11111111;
memory[6994]=8'b11111111;
memory[6995]=8'b11111111;
memory[6996]=8'b11111111;
memory[6997]=8'b11111111;
memory[6998]=8'b11111111;
memory[6999]=8'b11111111;
memory[7000]=8'b11111111;
memory[7001]=8'b11111111;
memory[7002]=8'b11111111;
memory[7003]=8'b11111111;
memory[7004]=8'b11111111;
memory[7005]=8'b11111111;
memory[7006]=8'b11111111;
memory[7007]=8'b11111111;
memory[7008]=8'b11111110;
memory[7009]=8'b00000111;
memory[7010]=8'b11111111;
memory[7011]=8'b11111111;
memory[7012]=8'b11111111;
memory[7013]=8'b11100001;
memory[7014]=8'b10011111;
memory[7015]=8'b11111111;
memory[7016]=8'b11111111;
memory[7017]=8'b11111111;
memory[7018]=8'b11111111;
memory[7019]=8'b11000000;
memory[7020]=8'b00000011;
memory[7021]=8'b11111111;
memory[7022]=8'b11111111;
memory[7023]=8'b11110000;
memory[7024]=8'b01111111;
memory[7025]=8'b11111111;
memory[7026]=8'b11111111;
memory[7027]=8'b11110010;
memory[7028]=8'b11111111;
memory[7029]=8'b11111111;
memory[7030]=8'b11111111;
memory[7031]=8'b11111111;
memory[7032]=8'b11111111;
memory[7033]=8'b11111111;
memory[7034]=8'b11111111;
memory[7035]=8'b11111111;
memory[7036]=8'b11111111;
memory[7037]=8'b11111111;
memory[7038]=8'b11111111;
memory[7039]=8'b11111111;
memory[7040]=8'b11111111;
memory[7041]=8'b11111111;
memory[7042]=8'b11111111;
memory[7043]=8'b11111111;
memory[7044]=8'b11111111;
memory[7045]=8'b11111111;
memory[7046]=8'b11111111;
memory[7047]=8'b11111111;
memory[7048]=8'b11111111;
memory[7049]=8'b11100000;
memory[7050]=8'b11111111;
memory[7051]=8'b11111111;
memory[7052]=8'b11111111;
memory[7053]=8'b11100001;
memory[7054]=8'b10011111;
memory[7055]=8'b11111111;
memory[7056]=8'b11111111;
memory[7057]=8'b11111111;
memory[7058]=8'b11111111;
memory[7059]=8'b11111100;
memory[7060]=8'b00000000;
memory[7061]=8'b00011111;
memory[7062]=8'b11100000;
memory[7063]=8'b00000011;
memory[7064]=8'b11111111;
memory[7065]=8'b11111111;
memory[7066]=8'b11111111;
memory[7067]=8'b11110000;
memory[7068]=8'b11111111;
memory[7069]=8'b11111111;
memory[7070]=8'b11111111;
memory[7071]=8'b11111111;
memory[7072]=8'b11111111;
memory[7073]=8'b11111111;
memory[7074]=8'b11111111;
memory[7075]=8'b11111111;
memory[7076]=8'b11111111;
memory[7077]=8'b11111111;
memory[7078]=8'b11111111;
memory[7079]=8'b11111111;
memory[7080]=8'b11111111;
memory[7081]=8'b11111111;
memory[7082]=8'b11111111;
memory[7083]=8'b11111111;
memory[7084]=8'b11111111;
memory[7085]=8'b11111111;
memory[7086]=8'b11111111;
memory[7087]=8'b11111111;
memory[7088]=8'b11111111;
memory[7089]=8'b11111000;
memory[7090]=8'b00011111;
memory[7091]=8'b11011111;
memory[7092]=8'b11111111;
memory[7093]=8'b11100001;
memory[7094]=8'b10001111;
memory[7095]=8'b11111111;
memory[7096]=8'b11111111;
memory[7097]=8'b11111111;
memory[7098]=8'b11111111;
memory[7099]=8'b11111111;
memory[7100]=8'b11000000;
memory[7101]=8'b00000000;
memory[7102]=8'b00000000;
memory[7103]=8'b00111111;
memory[7104]=8'b11111111;
memory[7105]=8'b11111111;
memory[7106]=8'b11111111;
memory[7107]=8'b11110000;
memory[7108]=8'b11111111;
memory[7109]=8'b11111111;
memory[7110]=8'b11111111;
memory[7111]=8'b11111111;
memory[7112]=8'b11111111;
memory[7113]=8'b11111111;
memory[7114]=8'b11111111;
memory[7115]=8'b11111111;
memory[7116]=8'b11111111;
memory[7117]=8'b11111111;
memory[7118]=8'b11111111;
memory[7119]=8'b11111111;
memory[7120]=8'b11111111;
memory[7121]=8'b11111111;
memory[7122]=8'b11111111;
memory[7123]=8'b11111111;
memory[7124]=8'b11111111;
memory[7125]=8'b11111111;
memory[7126]=8'b11111111;
memory[7127]=8'b11111111;
memory[7128]=8'b11111111;
memory[7129]=8'b11111111;
memory[7130]=8'b11000011;
memory[7131]=8'b11111111;
memory[7132]=8'b11111111;
memory[7133]=8'b11100001;
memory[7134]=8'b10001111;
memory[7135]=8'b11111111;
memory[7136]=8'b11111111;
memory[7137]=8'b11111111;
memory[7138]=8'b11111111;
memory[7139]=8'b11111111;
memory[7140]=8'b11111111;
memory[7141]=8'b11000000;
memory[7142]=8'b11111111;
memory[7143]=8'b11111111;
memory[7144]=8'b11111111;
memory[7145]=8'b11111111;
memory[7146]=8'b11111111;
memory[7147]=8'b11110000;
memory[7148]=8'b11111111;
memory[7149]=8'b11111111;
memory[7150]=8'b11111111;
memory[7151]=8'b11111111;
memory[7152]=8'b11111111;
memory[7153]=8'b11111111;
memory[7154]=8'b11111111;
memory[7155]=8'b11111111;
memory[7156]=8'b11111111;
memory[7157]=8'b11111111;
memory[7158]=8'b11111111;
memory[7159]=8'b11111111;
memory[7160]=8'b11111111;
memory[7161]=8'b11111111;
memory[7162]=8'b11111111;
memory[7163]=8'b11111111;
memory[7164]=8'b11111111;
memory[7165]=8'b11111111;
memory[7166]=8'b11111111;
memory[7167]=8'b11111111;
memory[7168]=8'b11111111;
memory[7169]=8'b11111111;
memory[7170]=8'b11111111;
memory[7171]=8'b11111111;
memory[7172]=8'b11111111;
memory[7173]=8'b11100001;
memory[7174]=8'b10001111;
memory[7175]=8'b11111111;
memory[7176]=8'b11111111;
memory[7177]=8'b11111111;
memory[7178]=8'b11111111;
memory[7179]=8'b11111111;
memory[7180]=8'b11111111;
memory[7181]=8'b11111111;
memory[7182]=8'b11111111;
memory[7183]=8'b11111111;
memory[7184]=8'b11111111;
memory[7185]=8'b11111111;
memory[7186]=8'b11111111;
memory[7187]=8'b11100000;
memory[7188]=8'b11111111;
memory[7189]=8'b11111111;
memory[7190]=8'b11111111;
memory[7191]=8'b11111111;
memory[7192]=8'b11111111;
memory[7193]=8'b11111111;
memory[7194]=8'b11111111;
memory[7195]=8'b11111111;
memory[7196]=8'b11111111;
memory[7197]=8'b11111111;
memory[7198]=8'b11111111;
memory[7199]=8'b11111111;
memory[7200]=8'b11111111;
memory[7201]=8'b11111111;
memory[7202]=8'b11111111;
memory[7203]=8'b11111111;
memory[7204]=8'b11111111;
memory[7205]=8'b11111111;
memory[7206]=8'b11111111;
memory[7207]=8'b11111111;
memory[7208]=8'b11111111;
memory[7209]=8'b11111111;
memory[7210]=8'b11111111;
memory[7211]=8'b11111111;
memory[7212]=8'b11111111;
memory[7213]=8'b11100011;
memory[7214]=8'b10001111;
memory[7215]=8'b11111111;
memory[7216]=8'b11111111;
memory[7217]=8'b11111111;
memory[7218]=8'b11111111;
memory[7219]=8'b11111111;
memory[7220]=8'b11111111;
memory[7221]=8'b11111111;
memory[7222]=8'b11111111;
memory[7223]=8'b11111111;
memory[7224]=8'b11111111;
memory[7225]=8'b11111111;
memory[7226]=8'b11111111;
memory[7227]=8'b11100100;
memory[7228]=8'b11111111;
memory[7229]=8'b11111111;
memory[7230]=8'b11111111;
memory[7231]=8'b11111111;
memory[7232]=8'b11111111;
memory[7233]=8'b11111111;
memory[7234]=8'b11111111;
memory[7235]=8'b11111111;
memory[7236]=8'b11111111;
memory[7237]=8'b11111111;
memory[7238]=8'b11111111;
memory[7239]=8'b11111111;
memory[7240]=8'b11111111;
memory[7241]=8'b11111111;
memory[7242]=8'b11111111;
memory[7243]=8'b11111111;
memory[7244]=8'b11111111;
memory[7245]=8'b11111111;
memory[7246]=8'b11111111;
memory[7247]=8'b11111111;
memory[7248]=8'b11111111;
memory[7249]=8'b11111111;
memory[7250]=8'b11111111;
memory[7251]=8'b11111111;
memory[7252]=8'b11111111;
memory[7253]=8'b11100001;
memory[7254]=8'b10000111;
memory[7255]=8'b11111111;
memory[7256]=8'b11111111;
memory[7257]=8'b11111111;
memory[7258]=8'b11111111;
memory[7259]=8'b11111111;
memory[7260]=8'b11111111;
memory[7261]=8'b11111111;
memory[7262]=8'b11111111;
memory[7263]=8'b11111111;
memory[7264]=8'b11111111;
memory[7265]=8'b11111111;
memory[7266]=8'b11111111;
memory[7267]=8'b11100100;
memory[7268]=8'b11111111;
memory[7269]=8'b11111111;
memory[7270]=8'b11111111;
memory[7271]=8'b11111111;
memory[7272]=8'b11111111;
memory[7273]=8'b11111111;
memory[7274]=8'b11111111;
memory[7275]=8'b11111111;
memory[7276]=8'b11111111;
memory[7277]=8'b11111111;
memory[7278]=8'b11111111;
memory[7279]=8'b11111111;
memory[7280]=8'b11111111;
memory[7281]=8'b11111111;
memory[7282]=8'b11111111;
memory[7283]=8'b11111111;
memory[7284]=8'b11111111;
memory[7285]=8'b11111111;
memory[7286]=8'b11111111;
memory[7287]=8'b11111111;
memory[7288]=8'b11111111;
memory[7289]=8'b11111111;
memory[7290]=8'b11111111;
memory[7291]=8'b11111111;
memory[7292]=8'b11111111;
memory[7293]=8'b11100001;
memory[7294]=8'b10000011;
memory[7295]=8'b11111111;
memory[7296]=8'b11111111;
memory[7297]=8'b11111111;
memory[7298]=8'b11111111;
memory[7299]=8'b11111111;
memory[7300]=8'b11111111;
memory[7301]=8'b11111111;
memory[7302]=8'b11111111;
memory[7303]=8'b11111111;
memory[7304]=8'b11111111;
memory[7305]=8'b11111111;
memory[7306]=8'b11111111;
memory[7307]=8'b11001100;
memory[7308]=8'b11111111;
memory[7309]=8'b11111111;
memory[7310]=8'b11111111;
memory[7311]=8'b11111111;
memory[7312]=8'b11111111;
memory[7313]=8'b11111111;
memory[7314]=8'b11111111;
memory[7315]=8'b11111111;
memory[7316]=8'b11111111;
memory[7317]=8'b11111111;
memory[7318]=8'b11111111;
memory[7319]=8'b11111111;
memory[7320]=8'b11111111;
memory[7321]=8'b11111111;
memory[7322]=8'b11111111;
memory[7323]=8'b11111111;
memory[7324]=8'b11111111;
memory[7325]=8'b11111111;
memory[7326]=8'b11111111;
memory[7327]=8'b11111111;
memory[7328]=8'b11111111;
memory[7329]=8'b11111111;
memory[7330]=8'b11111111;
memory[7331]=8'b11111111;
memory[7332]=8'b11111111;
memory[7333]=8'b11000000;
memory[7334]=8'b10000011;
memory[7335]=8'b11111111;
memory[7336]=8'b11111111;
memory[7337]=8'b11111111;
memory[7338]=8'b11111111;
memory[7339]=8'b11111111;
memory[7340]=8'b11111111;
memory[7341]=8'b11111111;
memory[7342]=8'b11111111;
memory[7343]=8'b11111111;
memory[7344]=8'b11111111;
memory[7345]=8'b11111111;
memory[7346]=8'b11111111;
memory[7347]=8'b11001100;
memory[7348]=8'b11111111;
memory[7349]=8'b11111111;
memory[7350]=8'b11111111;
memory[7351]=8'b11111111;
memory[7352]=8'b11111111;
memory[7353]=8'b11111111;
memory[7354]=8'b11111111;
memory[7355]=8'b11111111;
memory[7356]=8'b11111111;
memory[7357]=8'b11111111;
memory[7358]=8'b11111111;
memory[7359]=8'b11111111;
memory[7360]=8'b11111111;
memory[7361]=8'b11111111;
memory[7362]=8'b11111111;
memory[7363]=8'b11111111;
memory[7364]=8'b11111111;
memory[7365]=8'b11111111;
memory[7366]=8'b11111111;
memory[7367]=8'b11111111;
memory[7368]=8'b11111111;
memory[7369]=8'b11111111;
memory[7370]=8'b11111111;
memory[7371]=8'b11111111;
memory[7372]=8'b11111111;
memory[7373]=8'b11000000;
memory[7374]=8'b11000000;
memory[7375]=8'b11111111;
memory[7376]=8'b11111111;
memory[7377]=8'b11111111;
memory[7378]=8'b11111111;
memory[7379]=8'b11111111;
memory[7380]=8'b11111111;
memory[7381]=8'b11111111;
memory[7382]=8'b11111111;
memory[7383]=8'b11111111;
memory[7384]=8'b11111111;
memory[7385]=8'b11111111;
memory[7386]=8'b11111111;
memory[7387]=8'b11001100;
memory[7388]=8'b11111111;
memory[7389]=8'b11111111;
memory[7390]=8'b11111111;
memory[7391]=8'b11111111;
memory[7392]=8'b11111111;
memory[7393]=8'b11111111;
memory[7394]=8'b11111111;
memory[7395]=8'b11111111;
memory[7396]=8'b11111111;
memory[7397]=8'b11111111;
memory[7398]=8'b11111111;
memory[7399]=8'b11111111;
memory[7400]=8'b11111111;
memory[7401]=8'b11111111;
memory[7402]=8'b11111111;
memory[7403]=8'b11111111;
memory[7404]=8'b11111111;
memory[7405]=8'b11111111;
memory[7406]=8'b11111111;
memory[7407]=8'b11111111;
memory[7408]=8'b11111111;
memory[7409]=8'b11111111;
memory[7410]=8'b11111111;
memory[7411]=8'b11111111;
memory[7412]=8'b11111111;
memory[7413]=8'b10000000;
memory[7414]=8'b11000000;
memory[7415]=8'b00011111;
memory[7416]=8'b11111111;
memory[7417]=8'b11111111;
memory[7418]=8'b11111111;
memory[7419]=8'b11111111;
memory[7420]=8'b11111111;
memory[7421]=8'b11111111;
memory[7422]=8'b11111111;
memory[7423]=8'b11111111;
memory[7424]=8'b11111111;
memory[7425]=8'b11111111;
memory[7426]=8'b11111111;
memory[7427]=8'b10001100;
memory[7428]=8'b01111111;
memory[7429]=8'b11111111;
memory[7430]=8'b11111111;
memory[7431]=8'b11111111;
memory[7432]=8'b11111111;
memory[7433]=8'b11111111;
memory[7434]=8'b11111111;
memory[7435]=8'b11111111;
memory[7436]=8'b11111111;
memory[7437]=8'b11111111;
memory[7438]=8'b11111111;
memory[7439]=8'b11111111;
memory[7440]=8'b11111111;
memory[7441]=8'b11111111;
memory[7442]=8'b11111111;
memory[7443]=8'b11111111;
memory[7444]=8'b11111111;
memory[7445]=8'b11111111;
memory[7446]=8'b11111111;
memory[7447]=8'b11111111;
memory[7448]=8'b11111111;
memory[7449]=8'b11111111;
memory[7450]=8'b11111111;
memory[7451]=8'b11111111;
memory[7452]=8'b11111111;
memory[7453]=8'b00000000;
memory[7454]=8'b01100000;
memory[7455]=8'b00000011;
memory[7456]=8'b11111111;
memory[7457]=8'b11111111;
memory[7458]=8'b11111111;
memory[7459]=8'b11111111;
memory[7460]=8'b11111111;
memory[7461]=8'b11111111;
memory[7462]=8'b11111111;
memory[7463]=8'b11111111;
memory[7464]=8'b11111111;
memory[7465]=8'b11111111;
memory[7466]=8'b11111111;
memory[7467]=8'b00000000;
memory[7468]=8'b01111111;
memory[7469]=8'b11111111;
memory[7470]=8'b11111111;
memory[7471]=8'b11111111;
memory[7472]=8'b11111111;
memory[7473]=8'b11111111;
memory[7474]=8'b11111111;
memory[7475]=8'b11111111;
memory[7476]=8'b11111111;
memory[7477]=8'b11111111;
memory[7478]=8'b11111111;
memory[7479]=8'b11111111;
memory[7480]=8'b11111111;
memory[7481]=8'b11111111;
memory[7482]=8'b11111111;
memory[7483]=8'b11111111;
memory[7484]=8'b11111111;
memory[7485]=8'b11111111;
memory[7486]=8'b11111111;
memory[7487]=8'b11111111;
memory[7488]=8'b11111111;
memory[7489]=8'b11111111;
memory[7490]=8'b11111111;
memory[7491]=8'b11111111;
memory[7492]=8'b11111110;
memory[7493]=8'b00000000;
memory[7494]=8'b01100000;
memory[7495]=8'b00000000;
memory[7496]=8'b01111111;
memory[7497]=8'b11111111;
memory[7498]=8'b11111111;
memory[7499]=8'b11111111;
memory[7500]=8'b11111111;
memory[7501]=8'b11111111;
memory[7502]=8'b11111111;
memory[7503]=8'b11111111;
memory[7504]=8'b11111111;
memory[7505]=8'b11111111;
memory[7506]=8'b11111110;
memory[7507]=8'b00000000;
memory[7508]=8'b00111111;
memory[7509]=8'b11111111;
memory[7510]=8'b11111111;
memory[7511]=8'b11111111;
memory[7512]=8'b11111111;
memory[7513]=8'b11111111;
memory[7514]=8'b11111111;
memory[7515]=8'b11111111;
memory[7516]=8'b11111111;
memory[7517]=8'b11111111;
memory[7518]=8'b11111111;
memory[7519]=8'b11111111;
memory[7520]=8'b11111111;
memory[7521]=8'b11111111;
memory[7522]=8'b11111111;
memory[7523]=8'b11111111;
memory[7524]=8'b11111111;
memory[7525]=8'b11111111;
memory[7526]=8'b11111111;
memory[7527]=8'b11111111;
memory[7528]=8'b11111111;
memory[7529]=8'b11111111;
memory[7530]=8'b11111111;
memory[7531]=8'b11111111;
memory[7532]=8'b11111111;
memory[7533]=8'b11111111;
memory[7534]=8'b11110000;
memory[7535]=8'b00000000;
memory[7536]=8'b00000111;
memory[7537]=8'b11111111;
memory[7538]=8'b11111111;
memory[7539]=8'b11111111;
memory[7540]=8'b11111111;
memory[7541]=8'b11111111;
memory[7542]=8'b11111111;
memory[7543]=8'b11111111;
memory[7544]=8'b11111111;
memory[7545]=8'b11111111;
memory[7546]=8'b11110000;
memory[7547]=8'b00000000;
memory[7548]=8'b00011111;
memory[7549]=8'b11111111;
memory[7550]=8'b11111111;
memory[7551]=8'b11111111;
memory[7552]=8'b11111111;
memory[7553]=8'b11111111;
memory[7554]=8'b11111111;
memory[7555]=8'b11111111;
memory[7556]=8'b11111111;
memory[7557]=8'b11111111;
memory[7558]=8'b11111111;
memory[7559]=8'b11111111;
memory[7560]=8'b11111111;
memory[7561]=8'b11111111;
memory[7562]=8'b11111111;
memory[7563]=8'b11111111;
memory[7564]=8'b11111111;
memory[7565]=8'b11111111;
memory[7566]=8'b11111111;
memory[7567]=8'b11111111;
memory[7568]=8'b11111111;
memory[7569]=8'b11111111;
memory[7570]=8'b11111111;
memory[7571]=8'b11111111;
memory[7572]=8'b11111111;
memory[7573]=8'b11111111;
memory[7574]=8'b11110011;
memory[7575]=8'b11000000;
memory[7576]=8'b00000000;
memory[7577]=8'b11111111;
memory[7578]=8'b11111111;
memory[7579]=8'b11111111;
memory[7580]=8'b11111111;
memory[7581]=8'b11111111;
memory[7582]=8'b11111111;
memory[7583]=8'b11111111;
memory[7584]=8'b11111111;
memory[7585]=8'b11111111;
memory[7586]=8'b00000000;
memory[7587]=8'b00011000;
memory[7588]=8'b00011111;
memory[7589]=8'b11111111;
memory[7590]=8'b11111111;
memory[7591]=8'b11111111;
memory[7592]=8'b11111111;
memory[7593]=8'b11111111;
memory[7594]=8'b11111111;
memory[7595]=8'b11111111;
memory[7596]=8'b11111111;
memory[7597]=8'b11111111;
memory[7598]=8'b11111111;
memory[7599]=8'b11111111;
memory[7600]=8'b11111111;
memory[7601]=8'b11111111;
memory[7602]=8'b11111111;
memory[7603]=8'b11111111;
memory[7604]=8'b11111111;
memory[7605]=8'b11111111;
memory[7606]=8'b11111111;
memory[7607]=8'b11111111;
memory[7608]=8'b11111111;
memory[7609]=8'b11111111;
memory[7610]=8'b11111111;
memory[7611]=8'b11111111;
memory[7612]=8'b11111111;
memory[7613]=8'b11111111;
memory[7614]=8'b11111111;
memory[7615]=8'b11111111;
memory[7616]=8'b11111111;
memory[7617]=8'b11111111;
memory[7618]=8'b11111111;
memory[7619]=8'b11111111;
memory[7620]=8'b11111111;
memory[7621]=8'b11111111;
memory[7622]=8'b11111111;
memory[7623]=8'b11111111;
memory[7624]=8'b11111111;
memory[7625]=8'b11110000;
memory[7626]=8'b00000000;
memory[7627]=8'b00111111;
memory[7628]=8'b11111111;
memory[7629]=8'b11111111;
memory[7630]=8'b11111111;
memory[7631]=8'b11111111;
memory[7632]=8'b11111111;
memory[7633]=8'b11111111;
memory[7634]=8'b11111111;
memory[7635]=8'b11111111;
memory[7636]=8'b11111111;
memory[7637]=8'b11111111;
memory[7638]=8'b11111111;
memory[7639]=8'b11111111;
memory[7640]=8'b11111111;
memory[7641]=8'b11111111;
memory[7642]=8'b11111111;
memory[7643]=8'b11111111;
memory[7644]=8'b11111111;
memory[7645]=8'b11111111;
memory[7646]=8'b11111111;
memory[7647]=8'b11111111;
memory[7648]=8'b11111111;
memory[7649]=8'b11111111;
memory[7650]=8'b11111111;
memory[7651]=8'b11111111;
memory[7652]=8'b11111111;
memory[7653]=8'b11111111;
memory[7654]=8'b11111111;
memory[7655]=8'b11111111;
memory[7656]=8'b11111111;
memory[7657]=8'b11111111;
memory[7658]=8'b11111111;
memory[7659]=8'b11111111;
memory[7660]=8'b11111111;
memory[7661]=8'b11111111;
memory[7662]=8'b11111111;
memory[7663]=8'b11111111;
memory[7664]=8'b11111111;
memory[7665]=8'b11111111;
memory[7666]=8'b11111111;
memory[7667]=8'b11111111;
memory[7668]=8'b11111111;
memory[7669]=8'b11111111;
memory[7670]=8'b11111111;
memory[7671]=8'b11111111;
memory[7672]=8'b11111111;
memory[7673]=8'b11111111;
memory[7674]=8'b11111111;
memory[7675]=8'b11111111;
memory[7676]=8'b11111111;
memory[7677]=8'b11111111;
memory[7678]=8'b11111111;
memory[7679]=8'b11111111;
memory[7680]=8'b11111111;
memory[7681]=8'b11111111;
memory[7682]=8'b11111111;
memory[7683]=8'b11111111;
memory[7684]=8'b11111111;
memory[7685]=8'b11111111;
memory[7686]=8'b11111111;
memory[7687]=8'b11111111;
memory[7688]=8'b11111111;
memory[7689]=8'b11111111;
memory[7690]=8'b11111111;
memory[7691]=8'b11111111;
memory[7692]=8'b11111111;
memory[7693]=8'b11111111;
memory[7694]=8'b11111111;
memory[7695]=8'b11111111;
memory[7696]=8'b11111111;
memory[7697]=8'b11111111;
memory[7698]=8'b11111111;
memory[7699]=8'b11111111;
memory[7700]=8'b11111111;
memory[7701]=8'b11111111;
memory[7702]=8'b11111111;
memory[7703]=8'b11111111;
memory[7704]=8'b11111111;
memory[7705]=8'b11111111;
memory[7706]=8'b11111111;
memory[7707]=8'b11111111;
memory[7708]=8'b11111111;
memory[7709]=8'b11111111;
memory[7710]=8'b11111111;
memory[7711]=8'b11111111;
memory[7712]=8'b11111111;
memory[7713]=8'b11111111;
memory[7714]=8'b11111111;
memory[7715]=8'b11111111;
memory[7716]=8'b11111111;
memory[7717]=8'b11111111;
memory[7718]=8'b11111111;
memory[7719]=8'b11111111;
memory[7720]=8'b11111111;
memory[7721]=8'b11111111;
memory[7722]=8'b11111111;
memory[7723]=8'b11111111;
memory[7724]=8'b11111111;
memory[7725]=8'b11111111;
memory[7726]=8'b11111111;
memory[7727]=8'b11111111;
memory[7728]=8'b11111111;
memory[7729]=8'b11111111;
memory[7730]=8'b11111111;
memory[7731]=8'b11111111;
memory[7732]=8'b11111111;
memory[7733]=8'b11111111;
memory[7734]=8'b11111111;
memory[7735]=8'b11111111;
memory[7736]=8'b11111111;
memory[7737]=8'b11111111;
memory[7738]=8'b11111111;
memory[7739]=8'b11111111;
memory[7740]=8'b11111111;
memory[7741]=8'b11111111;
memory[7742]=8'b11111111;
memory[7743]=8'b11111111;
memory[7744]=8'b11111111;
memory[7745]=8'b11111111;
memory[7746]=8'b11111111;
memory[7747]=8'b11111111;
memory[7748]=8'b11111111;
memory[7749]=8'b11111111;
memory[7750]=8'b11111111;
memory[7751]=8'b11111111;
memory[7752]=8'b11111111;
memory[7753]=8'b11111111;
memory[7754]=8'b11111111;
memory[7755]=8'b11111111;
memory[7756]=8'b11111111;
memory[7757]=8'b11111111;
memory[7758]=8'b11111111;
memory[7759]=8'b11111111;
memory[7760]=8'b11111111;
memory[7761]=8'b11111111;
memory[7762]=8'b11111111;
memory[7763]=8'b11111111;
memory[7764]=8'b11111111;
memory[7765]=8'b11111111;
memory[7766]=8'b11111111;
memory[7767]=8'b11111111;
memory[7768]=8'b11111111;
memory[7769]=8'b11111111;
memory[7770]=8'b11111111;
memory[7771]=8'b11111111;
memory[7772]=8'b11111111;
memory[7773]=8'b11111111;
memory[7774]=8'b11111111;
memory[7775]=8'b11111111;
memory[7776]=8'b11111111;
memory[7777]=8'b11111111;
memory[7778]=8'b11111111;
memory[7779]=8'b11111111;
memory[7780]=8'b11111111;
memory[7781]=8'b11111111;
memory[7782]=8'b11111111;
memory[7783]=8'b11111111;
memory[7784]=8'b11111111;
memory[7785]=8'b11111111;
memory[7786]=8'b11111111;
memory[7787]=8'b11111111;
memory[7788]=8'b11111111;
memory[7789]=8'b11111111;
memory[7790]=8'b11111111;
memory[7791]=8'b11111111;
memory[7792]=8'b11111111;
memory[7793]=8'b11111111;
memory[7794]=8'b11111111;
memory[7795]=8'b11111111;
memory[7796]=8'b11111111;
memory[7797]=8'b11111111;
memory[7798]=8'b11111111;
memory[7799]=8'b11111111;
memory[7800]=8'b11111111;
memory[7801]=8'b11111111;
memory[7802]=8'b11111111;
memory[7803]=8'b11111111;
memory[7804]=8'b11111111;
memory[7805]=8'b11111111;
memory[7806]=8'b11111111;
memory[7807]=8'b11111111;
memory[7808]=8'b11111111;
memory[7809]=8'b11111111;
memory[7810]=8'b11111111;
memory[7811]=8'b11111111;
memory[7812]=8'b11111111;
memory[7813]=8'b11111111;
memory[7814]=8'b11111111;
memory[7815]=8'b11111111;
memory[7816]=8'b11111111;
memory[7817]=8'b11111111;
memory[7818]=8'b11111111;
memory[7819]=8'b11111111;
memory[7820]=8'b11111111;
memory[7821]=8'b11111111;
memory[7822]=8'b11111111;
memory[7823]=8'b11111111;
memory[7824]=8'b11111111;
memory[7825]=8'b11111111;
memory[7826]=8'b11111111;
memory[7827]=8'b11111111;
memory[7828]=8'b11111111;
memory[7829]=8'b11111111;
memory[7830]=8'b11111111;
memory[7831]=8'b11111111;
memory[7832]=8'b11111111;
memory[7833]=8'b11111111;
memory[7834]=8'b11111111;
memory[7835]=8'b11111111;
memory[7836]=8'b11111111;
memory[7837]=8'b11111111;
memory[7838]=8'b11111111;
memory[7839]=8'b11111111;
memory[7840]=8'b11111111;
memory[7841]=8'b11111111;
memory[7842]=8'b11111111;
memory[7843]=8'b11111111;
memory[7844]=8'b11111111;
memory[7845]=8'b11111111;
memory[7846]=8'b11111111;
memory[7847]=8'b11111111;
memory[7848]=8'b11111111;
memory[7849]=8'b11111111;
memory[7850]=8'b11111111;
memory[7851]=8'b11111111;
memory[7852]=8'b11111111;
memory[7853]=8'b11111111;
memory[7854]=8'b11111111;
memory[7855]=8'b11111111;
memory[7856]=8'b11111111;
memory[7857]=8'b11111111;
memory[7858]=8'b11111111;
memory[7859]=8'b11111111;
memory[7860]=8'b11111111;
memory[7861]=8'b11111111;
memory[7862]=8'b11111111;
memory[7863]=8'b11111111;
memory[7864]=8'b11111111;
memory[7865]=8'b11111111;
memory[7866]=8'b11111111;
memory[7867]=8'b11111111;
memory[7868]=8'b11111111;
memory[7869]=8'b11111111;
memory[7870]=8'b11111111;
memory[7871]=8'b11111111;
memory[7872]=8'b11111111;
memory[7873]=8'b11111111;
memory[7874]=8'b11111111;
memory[7875]=8'b11111111;
memory[7876]=8'b11111111;
memory[7877]=8'b11111111;
memory[7878]=8'b11111111;
memory[7879]=8'b11111111;
memory[7880]=8'b11111111;
memory[7881]=8'b11111111;
memory[7882]=8'b11111111;
memory[7883]=8'b11111111;
memory[7884]=8'b11111111;
memory[7885]=8'b11111111;
memory[7886]=8'b11111111;
memory[7887]=8'b11111111;
memory[7888]=8'b11111111;
memory[7889]=8'b11111111;
memory[7890]=8'b11111111;
memory[7891]=8'b11111111;
memory[7892]=8'b11111111;
memory[7893]=8'b11111111;
memory[7894]=8'b11111111;
memory[7895]=8'b11111111;
memory[7896]=8'b11111111;
memory[7897]=8'b11111111;
memory[7898]=8'b11111111;
memory[7899]=8'b11111111;
memory[7900]=8'b11111111;
memory[7901]=8'b11111111;
memory[7902]=8'b11111111;
memory[7903]=8'b11111111;
memory[7904]=8'b11111111;
memory[7905]=8'b11111111;
memory[7906]=8'b11111111;
memory[7907]=8'b11111111;
memory[7908]=8'b11111111;
memory[7909]=8'b11111111;
memory[7910]=8'b11111111;
memory[7911]=8'b11111111;
memory[7912]=8'b11111111;
memory[7913]=8'b11111111;
memory[7914]=8'b11111111;
memory[7915]=8'b11111111;
memory[7916]=8'b11111111;
memory[7917]=8'b11111111;
memory[7918]=8'b11111111;
memory[7919]=8'b11111111;
memory[7920]=8'b11111111;
memory[7921]=8'b11111111;
memory[7922]=8'b11111111;
memory[7923]=8'b11111111;
memory[7924]=8'b11111111;
memory[7925]=8'b11111111;
memory[7926]=8'b11111111;
memory[7927]=8'b11111111;
memory[7928]=8'b11111111;
memory[7929]=8'b11111111;
memory[7930]=8'b11111111;
memory[7931]=8'b11111111;
memory[7932]=8'b11111111;
memory[7933]=8'b11111111;
memory[7934]=8'b11111111;
memory[7935]=8'b11111111;
memory[7936]=8'b11111111;
memory[7937]=8'b11111111;
memory[7938]=8'b11111111;
memory[7939]=8'b11111111;
memory[7940]=8'b11111111;
memory[7941]=8'b11111111;
memory[7942]=8'b11111111;
memory[7943]=8'b11111111;
memory[7944]=8'b11111111;
memory[7945]=8'b11111111;
memory[7946]=8'b11111111;
memory[7947]=8'b11111111;
memory[7948]=8'b11111111;
memory[7949]=8'b11111111;
memory[7950]=8'b11111111;
memory[7951]=8'b11111111;
memory[7952]=8'b11111111;
memory[7953]=8'b11111111;
memory[7954]=8'b11111111;
memory[7955]=8'b11111111;
memory[7956]=8'b11111111;
memory[7957]=8'b11111111;
memory[7958]=8'b11111111;
memory[7959]=8'b11111111;
memory[7960]=8'b11111111;
memory[7961]=8'b11111111;
memory[7962]=8'b11111111;
memory[7963]=8'b11111111;
memory[7964]=8'b11111111;
memory[7965]=8'b11111111;
memory[7966]=8'b11111111;
memory[7967]=8'b11111111;
memory[7968]=8'b11111111;
memory[7969]=8'b11111111;
memory[7970]=8'b11111111;
memory[7971]=8'b11111111;
memory[7972]=8'b11111111;
memory[7973]=8'b11111111;
memory[7974]=8'b11111111;
memory[7975]=8'b11111111;
memory[7976]=8'b11111111;
memory[7977]=8'b11111111;
memory[7978]=8'b11111111;
memory[7979]=8'b11111111;
memory[7980]=8'b11111111;
memory[7981]=8'b11111111;
memory[7982]=8'b11111111;
memory[7983]=8'b11111111;
memory[7984]=8'b11111111;
memory[7985]=8'b11111111;
memory[7986]=8'b11111111;
memory[7987]=8'b11111111;
memory[7988]=8'b11111111;
memory[7989]=8'b11111111;
memory[7990]=8'b11111111;
memory[7991]=8'b11111111;
memory[7992]=8'b11111111;
memory[7993]=8'b11111111;
memory[7994]=8'b11111111;
memory[7995]=8'b11111111;
memory[7996]=8'b11111111;
memory[7997]=8'b11111111;
memory[7998]=8'b11111111;
memory[7999]=8'b11111111;

memory[8000]=8'b11111111;
memory[8001]=8'b11111111;
memory[8002]=8'b11111111;
memory[8003]=8'b11111111;
memory[8004]=8'b11111111;
memory[8005]=8'b11111111;
memory[8006]=8'b11111111;
memory[8007]=8'b11111111;
memory[8008]=8'b11111111;
memory[8009]=8'b11111111;
memory[8010]=8'b11111111;
memory[8011]=8'b11111111;
memory[8012]=8'b11111111;
memory[8013]=8'b11111111;
memory[8014]=8'b11111111;
memory[8015]=8'b11111111;
memory[8016]=8'b11111111;
memory[8017]=8'b11111111;
memory[8018]=8'b11111111;
memory[8019]=8'b11111111;
memory[8020]=8'b11111111;
memory[8021]=8'b11111111;
memory[8022]=8'b11111111;
memory[8023]=8'b11111111;
memory[8024]=8'b11111111;
memory[8025]=8'b11111111;
memory[8026]=8'b11111111;
memory[8027]=8'b11111111;
memory[8028]=8'b11111111;
memory[8029]=8'b11111111;
memory[8030]=8'b11111111;
memory[8031]=8'b11111111;
memory[8032]=8'b11111111;
memory[8033]=8'b11111111;
memory[8034]=8'b11111111;
memory[8035]=8'b11111111;
memory[8036]=8'b11111111;
memory[8037]=8'b11111111;
memory[8038]=8'b11111111;
memory[8039]=8'b11111111;
memory[8040]=8'b11111111;
memory[8041]=8'b11111111;
memory[8042]=8'b11111111;
memory[8043]=8'b11111111;
memory[8044]=8'b11111111;
memory[8045]=8'b11111111;
memory[8046]=8'b11111111;
memory[8047]=8'b11111111;
memory[8048]=8'b11111111;
memory[8049]=8'b11111111;
memory[8050]=8'b11111111;
memory[8051]=8'b11111111;
memory[8052]=8'b11111111;
memory[8053]=8'b11111111;
memory[8054]=8'b11111111;
memory[8055]=8'b11111111;
memory[8056]=8'b11111111;
memory[8057]=8'b11111111;
memory[8058]=8'b11111111;
memory[8059]=8'b11111111;
memory[8060]=8'b11111111;
memory[8061]=8'b11111111;
memory[8062]=8'b11111111;
memory[8063]=8'b11111111;
memory[8064]=8'b11111111;
memory[8065]=8'b11111111;
memory[8066]=8'b11111111;
memory[8067]=8'b11111111;
memory[8068]=8'b11111111;
memory[8069]=8'b11111111;
memory[8070]=8'b11111111;
memory[8071]=8'b11111111;
memory[8072]=8'b11111111;
memory[8073]=8'b11111111;
memory[8074]=8'b11111111;
memory[8075]=8'b11111111;
memory[8076]=8'b11111111;
memory[8077]=8'b11111111;
memory[8078]=8'b11111111;
memory[8079]=8'b11111111;
memory[8080]=8'b11111111;
memory[8081]=8'b11111111;
memory[8082]=8'b11111111;
memory[8083]=8'b11111111;
memory[8084]=8'b11111111;
memory[8085]=8'b11111111;
memory[8086]=8'b11111111;
memory[8087]=8'b11111111;
memory[8088]=8'b11111111;
memory[8089]=8'b11111111;
memory[8090]=8'b11111111;
memory[8091]=8'b11111111;
memory[8092]=8'b11111111;
memory[8093]=8'b11111111;
memory[8094]=8'b11111111;
memory[8095]=8'b11111111;
memory[8096]=8'b11111111;
memory[8097]=8'b11111111;
memory[8098]=8'b11111111;
memory[8099]=8'b11111111;
memory[8100]=8'b11111111;
memory[8101]=8'b11111111;
memory[8102]=8'b11111111;
memory[8103]=8'b11111111;
memory[8104]=8'b11111111;
memory[8105]=8'b11111111;
memory[8106]=8'b11111111;
memory[8107]=8'b11111111;
memory[8108]=8'b11111111;
memory[8109]=8'b11111111;
memory[8110]=8'b11111111;
memory[8111]=8'b11111111;
memory[8112]=8'b11111111;
memory[8113]=8'b11111111;
memory[8114]=8'b11111111;
memory[8115]=8'b11111111;
memory[8116]=8'b11111111;
memory[8117]=8'b11111111;
memory[8118]=8'b11111111;
memory[8119]=8'b11111111;
memory[8120]=8'b11111111;
memory[8121]=8'b11111111;
memory[8122]=8'b11111111;
memory[8123]=8'b11111111;
memory[8124]=8'b11111111;
memory[8125]=8'b11111111;
memory[8126]=8'b11111111;
memory[8127]=8'b11111111;
memory[8128]=8'b11111111;
memory[8129]=8'b11111111;
memory[8130]=8'b11111111;
memory[8131]=8'b11111111;
memory[8132]=8'b11111111;
memory[8133]=8'b11111111;
memory[8134]=8'b11111111;
memory[8135]=8'b11111111;
memory[8136]=8'b11111111;
memory[8137]=8'b11111111;
memory[8138]=8'b11111111;
memory[8139]=8'b11111111;
memory[8140]=8'b11111111;
memory[8141]=8'b11111111;
memory[8142]=8'b11111111;
memory[8143]=8'b11111111;
memory[8144]=8'b11111111;
memory[8145]=8'b11111111;
memory[8146]=8'b11111111;
memory[8147]=8'b11111111;
memory[8148]=8'b11111111;
memory[8149]=8'b11111111;
memory[8150]=8'b11111111;
memory[8151]=8'b11111111;
memory[8152]=8'b11111111;
memory[8153]=8'b11111111;
memory[8154]=8'b11111111;
memory[8155]=8'b11111111;
memory[8156]=8'b11111111;
memory[8157]=8'b11111111;
memory[8158]=8'b11111111;
memory[8159]=8'b11111111;
memory[8160]=8'b11111111;
memory[8161]=8'b11111111;
memory[8162]=8'b11111111;
memory[8163]=8'b11111111;
memory[8164]=8'b11111111;
memory[8165]=8'b11111111;
memory[8166]=8'b11111111;
memory[8167]=8'b11111111;
memory[8168]=8'b11111111;
memory[8169]=8'b11111111;
memory[8170]=8'b11111111;
memory[8171]=8'b11111111;
memory[8172]=8'b11111111;
memory[8173]=8'b11111111;
memory[8174]=8'b11111111;
memory[8175]=8'b11111111;
memory[8176]=8'b11111111;
memory[8177]=8'b11111111;
memory[8178]=8'b11111111;
memory[8179]=8'b11111111;
memory[8180]=8'b11111111;
memory[8181]=8'b11111111;
memory[8182]=8'b11111111;
memory[8183]=8'b11111111;
memory[8184]=8'b11111111;
memory[8185]=8'b11111111;
memory[8186]=8'b11111111;
memory[8187]=8'b11111111;
memory[8188]=8'b11111111;
memory[8189]=8'b11111111;
memory[8190]=8'b11111111;
memory[8191]=8'b11111111;
memory[8192]=8'b11111111;
memory[8193]=8'b11111111;
memory[8194]=8'b11111111;
memory[8195]=8'b11111111;
memory[8196]=8'b11111111;
memory[8197]=8'b11111111;
memory[8198]=8'b11111111;
memory[8199]=8'b11111111;
memory[8200]=8'b11111111;
memory[8201]=8'b11111111;
memory[8202]=8'b11111111;
memory[8203]=8'b11111111;
memory[8204]=8'b11111111;
memory[8205]=8'b11111111;
memory[8206]=8'b11111111;
memory[8207]=8'b11111111;
memory[8208]=8'b11111111;
memory[8209]=8'b11111111;
memory[8210]=8'b11111111;
memory[8211]=8'b11111111;
memory[8212]=8'b11111111;
memory[8213]=8'b11111111;
memory[8214]=8'b11111111;
memory[8215]=8'b11111111;
memory[8216]=8'b11111111;
memory[8217]=8'b11111111;
memory[8218]=8'b11111111;
memory[8219]=8'b11111111;
memory[8220]=8'b11111111;
memory[8221]=8'b11111111;
memory[8222]=8'b11111111;
memory[8223]=8'b11111111;
memory[8224]=8'b11111111;
memory[8225]=8'b11111111;
memory[8226]=8'b11111111;
memory[8227]=8'b11111111;
memory[8228]=8'b11111111;
memory[8229]=8'b11111111;
memory[8230]=8'b11111111;
memory[8231]=8'b11111111;
memory[8232]=8'b11111111;
memory[8233]=8'b11111111;
memory[8234]=8'b11111111;
memory[8235]=8'b11111111;
memory[8236]=8'b11111111;
memory[8237]=8'b11111111;
memory[8238]=8'b11111111;
memory[8239]=8'b11111111;
memory[8240]=8'b11111111;
memory[8241]=8'b11111111;
memory[8242]=8'b11111111;
memory[8243]=8'b11111111;
memory[8244]=8'b11111111;
memory[8245]=8'b11111111;
memory[8246]=8'b11111111;
memory[8247]=8'b11111111;
memory[8248]=8'b11111111;
memory[8249]=8'b11111111;
memory[8250]=8'b11111111;
memory[8251]=8'b11111111;
memory[8252]=8'b11111111;
memory[8253]=8'b11111111;
memory[8254]=8'b11111111;
memory[8255]=8'b11111111;
memory[8256]=8'b11111111;
memory[8257]=8'b11111111;
memory[8258]=8'b11111111;
memory[8259]=8'b11111111;
memory[8260]=8'b11111111;
memory[8261]=8'b11111111;
memory[8262]=8'b11111111;
memory[8263]=8'b11111111;
memory[8264]=8'b11111111;
memory[8265]=8'b11111111;
memory[8266]=8'b11111111;
memory[8267]=8'b11111111;
memory[8268]=8'b11111111;
memory[8269]=8'b11111111;
memory[8270]=8'b11111111;
memory[8271]=8'b11111111;
memory[8272]=8'b11111111;
memory[8273]=8'b11111111;
memory[8274]=8'b11111111;
memory[8275]=8'b11111111;
memory[8276]=8'b11111111;
memory[8277]=8'b11111111;
memory[8278]=8'b11111111;
memory[8279]=8'b11111111;
memory[8280]=8'b11111111;
memory[8281]=8'b11111111;
memory[8282]=8'b11111111;
memory[8283]=8'b11111111;
memory[8284]=8'b11111111;
memory[8285]=8'b11111111;
memory[8286]=8'b11111111;
memory[8287]=8'b11111111;
memory[8288]=8'b11111111;
memory[8289]=8'b11111111;
memory[8290]=8'b11111111;
memory[8291]=8'b11111111;
memory[8292]=8'b11111111;
memory[8293]=8'b11111111;
memory[8294]=8'b11111111;
memory[8295]=8'b11111111;
memory[8296]=8'b11111111;
memory[8297]=8'b11111111;
memory[8298]=8'b11111111;
memory[8299]=8'b11111111;
memory[8300]=8'b11111111;
memory[8301]=8'b11111111;
memory[8302]=8'b11111111;
memory[8303]=8'b11111111;
memory[8304]=8'b11111111;
memory[8305]=8'b11111111;
memory[8306]=8'b11111111;
memory[8307]=8'b11111111;
memory[8308]=8'b11111111;
memory[8309]=8'b11111111;
memory[8310]=8'b11111111;
memory[8311]=8'b11111111;
memory[8312]=8'b11111111;
memory[8313]=8'b11111111;
memory[8314]=8'b11111111;
memory[8315]=8'b11111111;
memory[8316]=8'b11111111;
memory[8317]=8'b11111111;
memory[8318]=8'b11111111;
memory[8319]=8'b11111111;
memory[8320]=8'b11111111;
memory[8321]=8'b11111111;
memory[8322]=8'b11111111;
memory[8323]=8'b11111111;
memory[8324]=8'b11111111;
memory[8325]=8'b11111111;
memory[8326]=8'b11111111;
memory[8327]=8'b11111111;
memory[8328]=8'b11111111;
memory[8329]=8'b11111111;
memory[8330]=8'b11111111;
memory[8331]=8'b11111111;
memory[8332]=8'b11111111;
memory[8333]=8'b11111111;
memory[8334]=8'b11111111;
memory[8335]=8'b11111111;
memory[8336]=8'b11111111;
memory[8337]=8'b11111111;
memory[8338]=8'b11111111;
memory[8339]=8'b11111111;
memory[8340]=8'b11111111;
memory[8341]=8'b11111111;
memory[8342]=8'b11111111;
memory[8343]=8'b11111111;
memory[8344]=8'b11111111;
memory[8345]=8'b11111111;
memory[8346]=8'b11111111;
memory[8347]=8'b11111111;
memory[8348]=8'b11111111;
memory[8349]=8'b11111111;
memory[8350]=8'b11111111;
memory[8351]=8'b11111111;
memory[8352]=8'b11111111;
memory[8353]=8'b11111111;
memory[8354]=8'b11111111;
memory[8355]=8'b11111111;
memory[8356]=8'b11111111;
memory[8357]=8'b11111111;
memory[8358]=8'b11111111;
memory[8359]=8'b11111111;
memory[8360]=8'b11111111;
memory[8361]=8'b11111111;
memory[8362]=8'b11111111;
memory[8363]=8'b11111111;
memory[8364]=8'b11111111;
memory[8365]=8'b11111111;
memory[8366]=8'b11111111;
memory[8367]=8'b11111111;
memory[8368]=8'b11111111;
memory[8369]=8'b11111111;
memory[8370]=8'b11111111;
memory[8371]=8'b11111111;
memory[8372]=8'b11111111;
memory[8373]=8'b11111111;
memory[8374]=8'b11111111;
memory[8375]=8'b11111111;
memory[8376]=8'b11111111;
memory[8377]=8'b11111111;
memory[8378]=8'b11111111;
memory[8379]=8'b11111111;
memory[8380]=8'b11111111;
memory[8381]=8'b11110000;
memory[8382]=8'b00011111;
memory[8383]=8'b11111111;
memory[8384]=8'b11111111;
memory[8385]=8'b11111111;
memory[8386]=8'b11111111;
memory[8387]=8'b11111111;
memory[8388]=8'b11111111;
memory[8389]=8'b11111111;
memory[8390]=8'b11111111;
memory[8391]=8'b11111111;
memory[8392]=8'b11111111;
memory[8393]=8'b11111111;
memory[8394]=8'b11111111;
memory[8395]=8'b11111111;
memory[8396]=8'b11111111;
memory[8397]=8'b11111111;
memory[8398]=8'b11111111;
memory[8399]=8'b11111111;
memory[8400]=8'b11111111;
memory[8401]=8'b11111111;
memory[8402]=8'b11111111;
memory[8403]=8'b11111111;
memory[8404]=8'b11111111;
memory[8405]=8'b11111111;
memory[8406]=8'b11111111;
memory[8407]=8'b11111111;
memory[8408]=8'b11111111;
memory[8409]=8'b11111111;
memory[8410]=8'b11111111;
memory[8411]=8'b11111111;
memory[8412]=8'b11111111;
memory[8413]=8'b11111111;
memory[8414]=8'b11111111;
memory[8415]=8'b11111111;
memory[8416]=8'b11111111;
memory[8417]=8'b11111111;
memory[8418]=8'b11111111;
memory[8419]=8'b11111111;
memory[8420]=8'b11111111;
memory[8421]=8'b00000000;
memory[8422]=8'b00000011;
memory[8423]=8'b11111111;
memory[8424]=8'b11111111;
memory[8425]=8'b11111111;
memory[8426]=8'b11111111;
memory[8427]=8'b11111111;
memory[8428]=8'b11111111;
memory[8429]=8'b11111111;
memory[8430]=8'b11111111;
memory[8431]=8'b11111111;
memory[8432]=8'b11111111;
memory[8433]=8'b11111111;
memory[8434]=8'b11111111;
memory[8435]=8'b11111111;
memory[8436]=8'b11111111;
memory[8437]=8'b11111111;
memory[8438]=8'b11111111;
memory[8439]=8'b11111111;
memory[8440]=8'b11111111;
memory[8441]=8'b11111111;
memory[8442]=8'b11111111;
memory[8443]=8'b11111111;
memory[8444]=8'b11111111;
memory[8445]=8'b11111111;
memory[8446]=8'b11111111;
memory[8447]=8'b11111111;
memory[8448]=8'b11111111;
memory[8449]=8'b11111111;
memory[8450]=8'b11111111;
memory[8451]=8'b11111111;
memory[8452]=8'b11111111;
memory[8453]=8'b11111111;
memory[8454]=8'b11111111;
memory[8455]=8'b11111111;
memory[8456]=8'b11111111;
memory[8457]=8'b11111111;
memory[8458]=8'b11111111;
memory[8459]=8'b11111111;
memory[8460]=8'b11111100;
memory[8461]=8'b00000000;
memory[8462]=8'b00000000;
memory[8463]=8'b11111111;
memory[8464]=8'b11111111;
memory[8465]=8'b11111111;
memory[8466]=8'b11111111;
memory[8467]=8'b11111111;
memory[8468]=8'b11111111;
memory[8469]=8'b11111111;
memory[8470]=8'b11111111;
memory[8471]=8'b11111111;
memory[8472]=8'b11111111;
memory[8473]=8'b11111111;
memory[8474]=8'b11111111;
memory[8475]=8'b11111111;
memory[8476]=8'b11111111;
memory[8477]=8'b11111111;
memory[8478]=8'b11111111;
memory[8479]=8'b11111111;
memory[8480]=8'b11111111;
memory[8481]=8'b11111111;
memory[8482]=8'b11111111;
memory[8483]=8'b11111111;
memory[8484]=8'b11111111;
memory[8485]=8'b11111111;
memory[8486]=8'b11111111;
memory[8487]=8'b11111111;
memory[8488]=8'b11111111;
memory[8489]=8'b11111111;
memory[8490]=8'b11111111;
memory[8491]=8'b11111111;
memory[8492]=8'b11111111;
memory[8493]=8'b11111111;
memory[8494]=8'b11111111;
memory[8495]=8'b11111111;
memory[8496]=8'b11111111;
memory[8497]=8'b11111111;
memory[8498]=8'b11111111;
memory[8499]=8'b11111111;
memory[8500]=8'b11111000;
memory[8501]=8'b00000000;
memory[8502]=8'b00000000;
memory[8503]=8'b01111111;
memory[8504]=8'b11111111;
memory[8505]=8'b11111111;
memory[8506]=8'b11111111;
memory[8507]=8'b11111111;
memory[8508]=8'b11111111;
memory[8509]=8'b11111111;
memory[8510]=8'b11111111;
memory[8511]=8'b11111111;
memory[8512]=8'b11111111;
memory[8513]=8'b11111111;
memory[8514]=8'b11111111;
memory[8515]=8'b11111111;
memory[8516]=8'b11111111;
memory[8517]=8'b11111111;
memory[8518]=8'b11111111;
memory[8519]=8'b11111111;
memory[8520]=8'b11111111;
memory[8521]=8'b11111111;
memory[8522]=8'b11111111;
memory[8523]=8'b11111111;
memory[8524]=8'b11111111;
memory[8525]=8'b11111111;
memory[8526]=8'b11111111;
memory[8527]=8'b11111111;
memory[8528]=8'b11111111;
memory[8529]=8'b11111111;
memory[8530]=8'b11111111;
memory[8531]=8'b11111111;
memory[8532]=8'b11111111;
memory[8533]=8'b11111111;
memory[8534]=8'b11111111;
memory[8535]=8'b11111111;
memory[8536]=8'b11111111;
memory[8537]=8'b11111111;
memory[8538]=8'b11111111;
memory[8539]=8'b11111111;
memory[8540]=8'b11110000;
memory[8541]=8'b00000000;
memory[8542]=8'b00000000;
memory[8543]=8'b00011111;
memory[8544]=8'b11111111;
memory[8545]=8'b11111111;
memory[8546]=8'b11111111;
memory[8547]=8'b11111111;
memory[8548]=8'b11111111;
memory[8549]=8'b11111111;
memory[8550]=8'b10011111;
memory[8551]=8'b11111111;
memory[8552]=8'b11111111;
memory[8553]=8'b11111111;
memory[8554]=8'b11111111;
memory[8555]=8'b11111111;
memory[8556]=8'b11111111;
memory[8557]=8'b11111111;
memory[8558]=8'b11111111;
memory[8559]=8'b11111111;
memory[8560]=8'b11111111;
memory[8561]=8'b11111111;
memory[8562]=8'b11111111;
memory[8563]=8'b11111111;
memory[8564]=8'b11111111;
memory[8565]=8'b11111111;
memory[8566]=8'b11111111;
memory[8567]=8'b11111111;
memory[8568]=8'b11111111;
memory[8569]=8'b11111111;
memory[8570]=8'b11111111;
memory[8571]=8'b11111111;
memory[8572]=8'b11111111;
memory[8573]=8'b11111111;
memory[8574]=8'b11111111;
memory[8575]=8'b11111111;
memory[8576]=8'b11111111;
memory[8577]=8'b11111111;
memory[8578]=8'b11111111;
memory[8579]=8'b11111111;
memory[8580]=8'b11100000;
memory[8581]=8'b00000000;
memory[8582]=8'b00000000;
memory[8583]=8'b00011111;
memory[8584]=8'b11111111;
memory[8585]=8'b11111111;
memory[8586]=8'b11111111;
memory[8587]=8'b11111111;
memory[8588]=8'b11111111;
memory[8589]=8'b11111111;
memory[8590]=8'b00001111;
memory[8591]=8'b11111111;
memory[8592]=8'b11111111;
memory[8593]=8'b11111111;
memory[8594]=8'b11111111;
memory[8595]=8'b11111111;
memory[8596]=8'b11111111;
memory[8597]=8'b11111111;
memory[8598]=8'b11111111;
memory[8599]=8'b11111111;
memory[8600]=8'b11111111;
memory[8601]=8'b11111111;
memory[8602]=8'b11111111;
memory[8603]=8'b11111111;
memory[8604]=8'b11111111;
memory[8605]=8'b11111111;
memory[8606]=8'b11111111;
memory[8607]=8'b11111111;
memory[8608]=8'b11111111;
memory[8609]=8'b11111111;
memory[8610]=8'b11111111;
memory[8611]=8'b11111111;
memory[8612]=8'b11111111;
memory[8613]=8'b11111111;
memory[8614]=8'b11111111;
memory[8615]=8'b11111111;
memory[8616]=8'b11111111;
memory[8617]=8'b11111111;
memory[8618]=8'b11111111;
memory[8619]=8'b11111111;
memory[8620]=8'b11100000;
memory[8621]=8'b00000000;
memory[8622]=8'b00000000;
memory[8623]=8'b00001111;
memory[8624]=8'b11111111;
memory[8625]=8'b11111111;
memory[8626]=8'b11111111;
memory[8627]=8'b11111111;
memory[8628]=8'b11111111;
memory[8629]=8'b11111111;
memory[8630]=8'b00001111;
memory[8631]=8'b11111111;
memory[8632]=8'b11111111;
memory[8633]=8'b11111111;
memory[8634]=8'b11111111;
memory[8635]=8'b11111111;
memory[8636]=8'b11111111;
memory[8637]=8'b11111111;
memory[8638]=8'b11111111;
memory[8639]=8'b11111111;
memory[8640]=8'b11111111;
memory[8641]=8'b11111111;
memory[8642]=8'b11111111;
memory[8643]=8'b11111111;
memory[8644]=8'b11111111;
memory[8645]=8'b11111111;
memory[8646]=8'b11111111;
memory[8647]=8'b11111111;
memory[8648]=8'b11111111;
memory[8649]=8'b11111111;
memory[8650]=8'b11111111;
memory[8651]=8'b11111111;
memory[8652]=8'b11111111;
memory[8653]=8'b11111111;
memory[8654]=8'b11111111;
memory[8655]=8'b11111111;
memory[8656]=8'b11111111;
memory[8657]=8'b11111111;
memory[8658]=8'b11111111;
memory[8659]=8'b11111111;
memory[8660]=8'b11100000;
memory[8661]=8'b00000000;
memory[8662]=8'b00000000;
memory[8663]=8'b00001111;
memory[8664]=8'b11111111;
memory[8665]=8'b11111111;
memory[8666]=8'b11111111;
memory[8667]=8'b11111111;
memory[8668]=8'b11111100;
memory[8669]=8'b11111111;
memory[8670]=8'b00000111;
memory[8671]=8'b11000000;
memory[8672]=8'b00111111;
memory[8673]=8'b11111111;
memory[8674]=8'b11111111;
memory[8675]=8'b11111111;
memory[8676]=8'b11111111;
memory[8677]=8'b11111111;
memory[8678]=8'b11111111;
memory[8679]=8'b11111111;
memory[8680]=8'b11111111;
memory[8681]=8'b11111111;
memory[8682]=8'b11111111;
memory[8683]=8'b11111111;
memory[8684]=8'b11111111;
memory[8685]=8'b11111111;
memory[8686]=8'b11111111;
memory[8687]=8'b11111111;
memory[8688]=8'b11111111;
memory[8689]=8'b11111111;
memory[8690]=8'b11111111;
memory[8691]=8'b11111111;
memory[8692]=8'b11111111;
memory[8693]=8'b11111111;
memory[8694]=8'b11111111;
memory[8695]=8'b11111111;
memory[8696]=8'b11111111;
memory[8697]=8'b11111111;
memory[8698]=8'b11111111;
memory[8699]=8'b11111111;
memory[8700]=8'b11100000;
memory[8701]=8'b00000000;
memory[8702]=8'b00000000;
memory[8703]=8'b00001111;
memory[8704]=8'b11111111;
memory[8705]=8'b11111111;
memory[8706]=8'b11111111;
memory[8707]=8'b11111111;
memory[8708]=8'b11110000;
memory[8709]=8'b00011111;
memory[8710]=8'b00001111;
memory[8711]=8'b00000001;
memory[8712]=8'b11111111;
memory[8713]=8'b11111111;
memory[8714]=8'b11111111;
memory[8715]=8'b11111111;
memory[8716]=8'b11111111;
memory[8717]=8'b11111111;
memory[8718]=8'b11111111;
memory[8719]=8'b11111111;
memory[8720]=8'b11111111;
memory[8721]=8'b11111111;
memory[8722]=8'b11111111;
memory[8723]=8'b11111111;
memory[8724]=8'b11111111;
memory[8725]=8'b11111111;
memory[8726]=8'b11111111;
memory[8727]=8'b11111111;
memory[8728]=8'b11111111;
memory[8729]=8'b11111111;
memory[8730]=8'b11111111;
memory[8731]=8'b11111111;
memory[8732]=8'b11111111;
memory[8733]=8'b11111111;
memory[8734]=8'b11111111;
memory[8735]=8'b11111111;
memory[8736]=8'b11111111;
memory[8737]=8'b11111111;
memory[8738]=8'b11111111;
memory[8739]=8'b11111111;
memory[8740]=8'b11100000;
memory[8741]=8'b00000000;
memory[8742]=8'b00000000;
memory[8743]=8'b00001111;
memory[8744]=8'b11111111;
memory[8745]=8'b11111111;
memory[8746]=8'b11111111;
memory[8747]=8'b11111111;
memory[8748]=8'b11111000;
memory[8749]=8'b00000111;
memory[8750]=8'b00001110;
memory[8751]=8'b00000011;
memory[8752]=8'b11111111;
memory[8753]=8'b11111111;
memory[8754]=8'b11111111;
memory[8755]=8'b11111111;
memory[8756]=8'b11111111;
memory[8757]=8'b11111111;
memory[8758]=8'b11111111;
memory[8759]=8'b11111111;
memory[8760]=8'b11111111;
memory[8761]=8'b11111111;
memory[8762]=8'b11111111;
memory[8763]=8'b11111111;
memory[8764]=8'b11111111;
memory[8765]=8'b11111111;
memory[8766]=8'b11111111;
memory[8767]=8'b11111111;
memory[8768]=8'b11111111;
memory[8769]=8'b11111111;
memory[8770]=8'b11111111;
memory[8771]=8'b11111111;
memory[8772]=8'b11111111;
memory[8773]=8'b11111111;
memory[8774]=8'b11111111;
memory[8775]=8'b11111111;
memory[8776]=8'b11111111;
memory[8777]=8'b11111111;
memory[8778]=8'b11111111;
memory[8779]=8'b11111111;
memory[8780]=8'b11110000;
memory[8781]=8'b00000000;
memory[8782]=8'b00000000;
memory[8783]=8'b00011111;
memory[8784]=8'b11111111;
memory[8785]=8'b11111111;
memory[8786]=8'b11111111;
memory[8787]=8'b11111111;
memory[8788]=8'b11111110;
memory[8789]=8'b00000001;
memory[8790]=8'b10001000;
memory[8791]=8'b00000000;
memory[8792]=8'b00011111;
memory[8793]=8'b11111111;
memory[8794]=8'b11111111;
memory[8795]=8'b11111111;
memory[8796]=8'b11111111;
memory[8797]=8'b11111111;
memory[8798]=8'b11111111;
memory[8799]=8'b11111111;
memory[8800]=8'b11111111;
memory[8801]=8'b11111111;
memory[8802]=8'b11111111;
memory[8803]=8'b11111111;
memory[8804]=8'b11111111;
memory[8805]=8'b11111111;
memory[8806]=8'b11111111;
memory[8807]=8'b11111111;
memory[8808]=8'b11111111;
memory[8809]=8'b11111111;
memory[8810]=8'b11111111;
memory[8811]=8'b11111111;
memory[8812]=8'b11111111;
memory[8813]=8'b11111111;
memory[8814]=8'b11111111;
memory[8815]=8'b11111111;
memory[8816]=8'b11111111;
memory[8817]=8'b11111111;
memory[8818]=8'b11111111;
memory[8819]=8'b11111111;
memory[8820]=8'b11110000;
memory[8821]=8'b00000000;
memory[8822]=8'b00000000;
memory[8823]=8'b00111111;
memory[8824]=8'b11111111;
memory[8825]=8'b11111111;
memory[8826]=8'b11111111;
memory[8827]=8'b11111111;
memory[8828]=8'b11111111;
memory[8829]=8'b11111000;
memory[8830]=8'b11001000;
memory[8831]=8'b00000011;
memory[8832]=8'b11111111;
memory[8833]=8'b11111111;
memory[8834]=8'b11111111;
memory[8835]=8'b11111111;
memory[8836]=8'b11111111;
memory[8837]=8'b11111111;
memory[8838]=8'b11111111;
memory[8839]=8'b11111111;
memory[8840]=8'b11111111;
memory[8841]=8'b11111111;
memory[8842]=8'b11111111;
memory[8843]=8'b11111111;
memory[8844]=8'b11111111;
memory[8845]=8'b11111111;
memory[8846]=8'b11111111;
memory[8847]=8'b11111111;
memory[8848]=8'b11111111;
memory[8849]=8'b11111111;
memory[8850]=8'b11111111;
memory[8851]=8'b11111111;
memory[8852]=8'b11111111;
memory[8853]=8'b11111111;
memory[8854]=8'b11111111;
memory[8855]=8'b11111111;
memory[8856]=8'b11111111;
memory[8857]=8'b11111111;
memory[8858]=8'b11111111;
memory[8859]=8'b11111111;
memory[8860]=8'b11111000;
memory[8861]=8'b00000000;
memory[8862]=8'b00000000;
memory[8863]=8'b01111111;
memory[8864]=8'b11111111;
memory[8865]=8'b11111111;
memory[8866]=8'b11111111;
memory[8867]=8'b11111111;
memory[8868]=8'b11100000;
memory[8869]=8'b00111110;
memory[8870]=8'b01001000;
memory[8871]=8'b00111111;
memory[8872]=8'b11111111;
memory[8873]=8'b11111111;
memory[8874]=8'b11111111;
memory[8875]=8'b11111111;
memory[8876]=8'b11111111;
memory[8877]=8'b11111111;
memory[8878]=8'b11111111;
memory[8879]=8'b11111111;
memory[8880]=8'b11111111;
memory[8881]=8'b11111111;
memory[8882]=8'b11111111;
memory[8883]=8'b11111111;
memory[8884]=8'b11111111;
memory[8885]=8'b11111111;
memory[8886]=8'b11111111;
memory[8887]=8'b11111111;
memory[8888]=8'b11111111;
memory[8889]=8'b11111111;
memory[8890]=8'b11111111;
memory[8891]=8'b11111111;
memory[8892]=8'b11111111;
memory[8893]=8'b11111111;
memory[8894]=8'b11111111;
memory[8895]=8'b11111111;
memory[8896]=8'b11111111;
memory[8897]=8'b11111111;
memory[8898]=8'b11111111;
memory[8899]=8'b11111111;
memory[8900]=8'b11111110;
memory[8901]=8'b00000000;
memory[8902]=8'b00000000;
memory[8903]=8'b11111111;
memory[8904]=8'b11111111;
memory[8905]=8'b11111111;
memory[8906]=8'b11111111;
memory[8907]=8'b11111111;
memory[8908]=8'b00000000;
memory[8909]=8'b00000001;
memory[8910]=8'b11111111;
memory[8911]=8'b11100000;
memory[8912]=8'b00001111;
memory[8913]=8'b11111111;
memory[8914]=8'b11111111;
memory[8915]=8'b11111111;
memory[8916]=8'b11111111;
memory[8917]=8'b11111111;
memory[8918]=8'b11111111;
memory[8919]=8'b11111111;
memory[8920]=8'b11111111;
memory[8921]=8'b11111111;
memory[8922]=8'b11111111;
memory[8923]=8'b11111111;
memory[8924]=8'b11111111;
memory[8925]=8'b11111111;
memory[8926]=8'b11111111;
memory[8927]=8'b11111111;
memory[8928]=8'b11111111;
memory[8929]=8'b11111111;
memory[8930]=8'b11111111;
memory[8931]=8'b11111111;
memory[8932]=8'b11111111;
memory[8933]=8'b11111111;
memory[8934]=8'b11111111;
memory[8935]=8'b11111111;
memory[8936]=8'b11111111;
memory[8937]=8'b11111111;
memory[8938]=8'b11111111;
memory[8939]=8'b11111111;
memory[8940]=8'b11111111;
memory[8941]=8'b10000000;
memory[8942]=8'b00000011;
memory[8943]=8'b11111111;
memory[8944]=8'b11111111;
memory[8945]=8'b11111111;
memory[8946]=8'b11111111;
memory[8947]=8'b11111100;
memory[8948]=8'b00000000;
memory[8949]=8'b00011100;
memory[8950]=8'b11111111;
memory[8951]=8'b00000000;
memory[8952]=8'b00000011;
memory[8953]=8'b11111111;
memory[8954]=8'b11111111;
memory[8955]=8'b11111111;
memory[8956]=8'b11111111;
memory[8957]=8'b11111111;
memory[8958]=8'b11111111;
memory[8959]=8'b11111111;
memory[8960]=8'b11111111;
memory[8961]=8'b11111111;
memory[8962]=8'b11111111;
memory[8963]=8'b11111111;
memory[8964]=8'b11111111;
memory[8965]=8'b11111111;
memory[8966]=8'b11111111;
memory[8967]=8'b11111111;
memory[8968]=8'b11111111;
memory[8969]=8'b11111111;
memory[8970]=8'b11111111;
memory[8971]=8'b11111111;
memory[8972]=8'b11111111;
memory[8973]=8'b11111111;
memory[8974]=8'b11111111;
memory[8975]=8'b11111111;
memory[8976]=8'b11111111;
memory[8977]=8'b11111111;
memory[8978]=8'b11111111;
memory[8979]=8'b11111111;
memory[8980]=8'b11111111;
memory[8981]=8'b11111000;
memory[8982]=8'b00111111;
memory[8983]=8'b11111111;
memory[8984]=8'b11111111;
memory[8985]=8'b11110011;
memory[8986]=8'b11111111;
memory[8987]=8'b11111111;
memory[8988]=8'b11111110;
memory[8989]=8'b00000000;
memory[8990]=8'b00111111;
memory[8991]=8'b01100011;
memory[8992]=8'b11111111;
memory[8993]=8'b11111111;
memory[8994]=8'b11111111;
memory[8995]=8'b11111111;
memory[8996]=8'b11111111;
memory[8997]=8'b11111111;
memory[8998]=8'b11111111;
memory[8999]=8'b11111111;
memory[9000]=8'b11111111;
memory[9001]=8'b11111111;
memory[9002]=8'b11111111;
memory[9003]=8'b11111111;
memory[9004]=8'b11111111;
memory[9005]=8'b11111111;
memory[9006]=8'b11111111;
memory[9007]=8'b11111111;
memory[9008]=8'b11111111;
memory[9009]=8'b11111111;
memory[9010]=8'b11111111;
memory[9011]=8'b11111111;
memory[9012]=8'b11111111;
memory[9013]=8'b11111111;
memory[9014]=8'b11111111;
memory[9015]=8'b11111111;
memory[9016]=8'b11111111;
memory[9017]=8'b11111111;
memory[9018]=8'b11111111;
memory[9019]=8'b11111111;
memory[9020]=8'b11111111;
memory[9021]=8'b11111111;
memory[9022]=8'b11111111;
memory[9023]=8'b11111111;
memory[9024]=8'b11111111;
memory[9025]=8'b00000111;
memory[9026]=8'b11111111;
memory[9027]=8'b11111111;
memory[9028]=8'b11110000;
memory[9029]=8'b00000000;
memory[9030]=8'b00000000;
memory[9031]=8'b00000011;
memory[9032]=8'b11111111;
memory[9033]=8'b11111111;
memory[9034]=8'b11111111;
memory[9035]=8'b11111111;
memory[9036]=8'b11111111;
memory[9037]=8'b11111111;
memory[9038]=8'b11111111;
memory[9039]=8'b11111111;
memory[9040]=8'b11111111;
memory[9041]=8'b11111111;
memory[9042]=8'b11111111;
memory[9043]=8'b11111111;
memory[9044]=8'b11111111;
memory[9045]=8'b11111111;
memory[9046]=8'b11111111;
memory[9047]=8'b11111111;
memory[9048]=8'b11111111;
memory[9049]=8'b11111111;
memory[9050]=8'b11111111;
memory[9051]=8'b11111111;
memory[9052]=8'b11111111;
memory[9053]=8'b11111111;
memory[9054]=8'b11111111;
memory[9055]=8'b11111111;
memory[9056]=8'b11111111;
memory[9057]=8'b11111111;
memory[9058]=8'b11111111;
memory[9059]=8'b11111111;
memory[9060]=8'b11111111;
memory[9061]=8'b11111111;
memory[9062]=8'b11111111;
memory[9063]=8'b11111111;
memory[9064]=8'b11111100;
memory[9065]=8'b00001111;
memory[9066]=8'b11111111;
memory[9067]=8'b11111111;
memory[9068]=8'b11000001;
memory[9069]=8'b00000010;
memory[9070]=8'b00000011;
memory[9071]=8'b00000001;
memory[9072]=8'b11111111;
memory[9073]=8'b11111111;
memory[9074]=8'b11111111;
memory[9075]=8'b11111111;
memory[9076]=8'b11111111;
memory[9077]=8'b11111111;
memory[9078]=8'b11111111;
memory[9079]=8'b11111111;
memory[9080]=8'b11111111;
memory[9081]=8'b11111111;
memory[9082]=8'b11111111;
memory[9083]=8'b11111111;
memory[9084]=8'b11111111;
memory[9085]=8'b11111111;
memory[9086]=8'b11111111;
memory[9087]=8'b11111111;
memory[9088]=8'b11111111;
memory[9089]=8'b11111111;
memory[9090]=8'b11111111;
memory[9091]=8'b11111111;
memory[9092]=8'b11111111;
memory[9093]=8'b11111111;
memory[9094]=8'b11111111;
memory[9095]=8'b11111111;
memory[9096]=8'b11111111;
memory[9097]=8'b11111111;
memory[9098]=8'b11111111;
memory[9099]=8'b11111111;
memory[9100]=8'b11111111;
memory[9101]=8'b11111111;
memory[9102]=8'b11111111;
memory[9103]=8'b11111111;
memory[9104]=8'b11111000;
memory[9105]=8'b00111100;
memory[9106]=8'b00000001;
memory[9107]=8'b11111111;
memory[9108]=8'b00011111;
memory[9109]=8'b10000000;
memory[9110]=8'b00000011;
memory[9111]=8'b00000000;
memory[9112]=8'b00111111;
memory[9113]=8'b11111111;
memory[9114]=8'b11111111;
memory[9115]=8'b11111111;
memory[9116]=8'b11111111;
memory[9117]=8'b11111111;
memory[9118]=8'b11111111;
memory[9119]=8'b11111111;
memory[9120]=8'b11111111;
memory[9121]=8'b11111111;
memory[9122]=8'b11111111;
memory[9123]=8'b11111111;
memory[9124]=8'b11111111;
memory[9125]=8'b11111111;
memory[9126]=8'b11111111;
memory[9127]=8'b11111111;
memory[9128]=8'b11111111;
memory[9129]=8'b11111111;
memory[9130]=8'b11111111;
memory[9131]=8'b11111111;
memory[9132]=8'b11111111;
memory[9133]=8'b11111111;
memory[9134]=8'b11111111;
memory[9135]=8'b11111111;
memory[9136]=8'b11111111;
memory[9137]=8'b11111111;
memory[9138]=8'b11111111;
memory[9139]=8'b11111111;
memory[9140]=8'b11111111;
memory[9141]=8'b11111111;
memory[9142]=8'b11111111;
memory[9143]=8'b11111111;
memory[9144]=8'b11111000;
memory[9145]=8'b00110000;
memory[9146]=8'b00000000;
memory[9147]=8'b01111111;
memory[9148]=8'b11111111;
memory[9149]=8'b00000011;
memory[9150]=8'b00000001;
memory[9151]=8'b10000000;
memory[9152]=8'b00011111;
memory[9153]=8'b11111111;
memory[9154]=8'b11111111;
memory[9155]=8'b11111111;
memory[9156]=8'b11111111;
memory[9157]=8'b11111111;
memory[9158]=8'b11111111;
memory[9159]=8'b11111111;
memory[9160]=8'b11111111;
memory[9161]=8'b11111111;
memory[9162]=8'b11111111;
memory[9163]=8'b11111111;
memory[9164]=8'b11111111;
memory[9165]=8'b11111111;
memory[9166]=8'b11111111;
memory[9167]=8'b11111111;
memory[9168]=8'b11111111;
memory[9169]=8'b11111111;
memory[9170]=8'b11111111;
memory[9171]=8'b11111111;
memory[9172]=8'b11111111;
memory[9173]=8'b11111111;
memory[9174]=8'b11111111;
memory[9175]=8'b11111111;
memory[9176]=8'b11111111;
memory[9177]=8'b11111111;
memory[9178]=8'b11111111;
memory[9179]=8'b11111111;
memory[9180]=8'b11111111;
memory[9181]=8'b11111111;
memory[9182]=8'b11111111;
memory[9183]=8'b11111111;
memory[9184]=8'b11111100;
memory[9185]=8'b01100000;
memory[9186]=8'b11111110;
memory[9187]=8'b00011111;
memory[9188]=8'b11111100;
memory[9189]=8'b00000111;
memory[9190]=8'b00000001;
memory[9191]=8'b10000000;
memory[9192]=8'b00001111;
memory[9193]=8'b11111111;
memory[9194]=8'b11111111;
memory[9195]=8'b11111111;
memory[9196]=8'b11111111;
memory[9197]=8'b11111111;
memory[9198]=8'b11111111;
memory[9199]=8'b11111111;
memory[9200]=8'b11111111;
memory[9201]=8'b11111111;
memory[9202]=8'b11111111;
memory[9203]=8'b11111111;
memory[9204]=8'b11111111;
memory[9205]=8'b11111111;
memory[9206]=8'b11111111;
memory[9207]=8'b11111111;
memory[9208]=8'b11111111;
memory[9209]=8'b11111111;
memory[9210]=8'b11111111;
memory[9211]=8'b11111111;
memory[9212]=8'b11111111;
memory[9213]=8'b11111111;
memory[9214]=8'b11111111;
memory[9215]=8'b11111111;
memory[9216]=8'b11111111;
memory[9217]=8'b11111111;
memory[9218]=8'b11111111;
memory[9219]=8'b11111111;
memory[9220]=8'b11111111;
memory[9221]=8'b11111111;
memory[9222]=8'b11111111;
memory[9223]=8'b11111100;
memory[9224]=8'b00001110;
memory[9225]=8'b01101111;
memory[9226]=8'b10011000;
memory[9227]=8'b11111111;
memory[9228]=8'b11111100;
memory[9229]=8'b00001100;
memory[9230]=8'b11100001;
memory[9231]=8'b10000010;
memory[9232]=8'b00001111;
memory[9233]=8'b11111111;
memory[9234]=8'b11111111;
memory[9235]=8'b11111111;
memory[9236]=8'b11111111;
memory[9237]=8'b11111111;
memory[9238]=8'b11111111;
memory[9239]=8'b11111111;
memory[9240]=8'b11111111;
memory[9241]=8'b11111111;
memory[9242]=8'b11111111;
memory[9243]=8'b11111111;
memory[9244]=8'b11111111;
memory[9245]=8'b11111111;
memory[9246]=8'b11111111;
memory[9247]=8'b11111111;
memory[9248]=8'b11111111;
memory[9249]=8'b11111111;
memory[9250]=8'b11111111;
memory[9251]=8'b11111111;
memory[9252]=8'b11111111;
memory[9253]=8'b11111111;
memory[9254]=8'b11111111;
memory[9255]=8'b11111111;
memory[9256]=8'b11111111;
memory[9257]=8'b11111111;
memory[9258]=8'b11111111;
memory[9259]=8'b11111111;
memory[9260]=8'b11111111;
memory[9261]=8'b11111111;
memory[9262]=8'b11111111;
memory[9263]=8'b11100000;
memory[9264]=8'b00000011;
memory[9265]=8'b01100000;
memory[9266]=8'b00000000;
memory[9267]=8'b00111111;
memory[9268]=8'b11111100;
memory[9269]=8'b01111000;
memory[9270]=8'b11100000;
memory[9271]=8'b10000011;
memory[9272]=8'b10000111;
memory[9273]=8'b11111111;
memory[9274]=8'b11111111;
memory[9275]=8'b11111111;
memory[9276]=8'b11111111;
memory[9277]=8'b11111111;
memory[9278]=8'b11111111;
memory[9279]=8'b11111111;
memory[9280]=8'b11111111;
memory[9281]=8'b11111111;
memory[9282]=8'b11111111;
memory[9283]=8'b11111111;
memory[9284]=8'b11111111;
memory[9285]=8'b11111111;
memory[9286]=8'b11111111;
memory[9287]=8'b11111111;
memory[9288]=8'b11111111;
memory[9289]=8'b11111111;
memory[9290]=8'b11111111;
memory[9291]=8'b11111111;
memory[9292]=8'b11111111;
memory[9293]=8'b11111111;
memory[9294]=8'b11111111;
memory[9295]=8'b11111111;
memory[9296]=8'b11111111;
memory[9297]=8'b11111111;
memory[9298]=8'b11111111;
memory[9299]=8'b11111111;
memory[9300]=8'b11111111;
memory[9301]=8'b11111111;
memory[9302]=8'b11111111;
memory[9303]=8'b11000000;
memory[9304]=8'b00111111;
memory[9305]=8'b11110000;
memory[9306]=8'b00000000;
memory[9307]=8'b00001111;
memory[9308]=8'b11111111;
memory[9309]=8'b11111001;
memory[9310]=8'b11110000;
memory[9311]=8'b11000001;
memory[9312]=8'b11110011;
memory[9313]=8'b11111111;
memory[9314]=8'b11111111;
memory[9315]=8'b11111111;
memory[9316]=8'b11111111;
memory[9317]=8'b11111111;
memory[9318]=8'b11111111;
memory[9319]=8'b11111111;
memory[9320]=8'b11111111;
memory[9321]=8'b11111111;
memory[9322]=8'b11111111;
memory[9323]=8'b11111111;
memory[9324]=8'b11111111;
memory[9325]=8'b11111111;
memory[9326]=8'b11111111;
memory[9327]=8'b11111111;
memory[9328]=8'b11111111;
memory[9329]=8'b11111111;
memory[9330]=8'b11111111;
memory[9331]=8'b11111111;
memory[9332]=8'b11111111;
memory[9333]=8'b11111111;
memory[9334]=8'b11111111;
memory[9335]=8'b11111111;
memory[9336]=8'b11111111;
memory[9337]=8'b11111111;
memory[9338]=8'b11111111;
memory[9339]=8'b11111111;
memory[9340]=8'b11111111;
memory[9341]=8'b11111111;
memory[9342]=8'b11111111;
memory[9343]=8'b10000001;
memory[9344]=8'b11111111;
memory[9345]=8'b11111111;
memory[9346]=8'b00000000;
memory[9347]=8'b00000111;
memory[9348]=8'b11111111;
memory[9349]=8'b11110011;
memory[9350]=8'b11111000;
memory[9351]=8'b11100001;
memory[9352]=8'b11111111;
memory[9353]=8'b11111111;
memory[9354]=8'b11111111;
memory[9355]=8'b11111111;
memory[9356]=8'b11111111;
memory[9357]=8'b11111111;
memory[9358]=8'b11111111;
memory[9359]=8'b11111111;
memory[9360]=8'b11111111;
memory[9361]=8'b11111111;
memory[9362]=8'b11111111;
memory[9363]=8'b11111111;
memory[9364]=8'b11111111;
memory[9365]=8'b11111111;
memory[9366]=8'b11111111;
memory[9367]=8'b11111111;
memory[9368]=8'b11111111;
memory[9369]=8'b11111111;
memory[9370]=8'b11111111;
memory[9371]=8'b11111111;
memory[9372]=8'b11111111;
memory[9373]=8'b11111111;
memory[9374]=8'b11111111;
memory[9375]=8'b11111111;
memory[9376]=8'b11111111;
memory[9377]=8'b11111111;
memory[9378]=8'b11111111;
memory[9379]=8'b11111111;
memory[9380]=8'b11111111;
memory[9381]=8'b11111111;
memory[9382]=8'b11111111;
memory[9383]=8'b00001111;
memory[9384]=8'b10000011;
memory[9385]=8'b10000000;
memory[9386]=8'b11000000;
memory[9387]=8'b00000011;
memory[9388]=8'b11111111;
memory[9389]=8'b11100011;
memory[9390]=8'b11111000;
memory[9391]=8'b11110001;
memory[9392]=8'b11111111;
memory[9393]=8'b11111111;
memory[9394]=8'b11111111;
memory[9395]=8'b11111111;
memory[9396]=8'b11111111;
memory[9397]=8'b11111111;
memory[9398]=8'b11111111;
memory[9399]=8'b11111111;
memory[9400]=8'b11111111;
memory[9401]=8'b11111111;
memory[9402]=8'b11111111;
memory[9403]=8'b11111111;
memory[9404]=8'b11111111;
memory[9405]=8'b11111111;
memory[9406]=8'b11111111;
memory[9407]=8'b11111111;
memory[9408]=8'b11111111;
memory[9409]=8'b11111111;
memory[9410]=8'b11111111;
memory[9411]=8'b11111111;
memory[9412]=8'b11111111;
memory[9413]=8'b11111111;
memory[9414]=8'b11111111;
memory[9415]=8'b11111111;
memory[9416]=8'b11111111;
memory[9417]=8'b11111111;
memory[9418]=8'b11000000;
memory[9419]=8'b00000001;
memory[9420]=8'b11111111;
memory[9421]=8'b11111111;
memory[9422]=8'b11111110;
memory[9423]=8'b00001100;
memory[9424]=8'b00000111;
memory[9425]=8'b10000000;
memory[9426]=8'b01110000;
memory[9427]=8'b01111001;
memory[9428]=8'b11111111;
memory[9429]=8'b11100111;
memory[9430]=8'b11111000;
memory[9431]=8'b11111101;
memory[9432]=8'b11111111;
memory[9433]=8'b11111111;
memory[9434]=8'b11111111;
memory[9435]=8'b11111111;
memory[9436]=8'b11111111;
memory[9437]=8'b11111111;
memory[9438]=8'b11111111;
memory[9439]=8'b11111111;
memory[9440]=8'b11111111;
memory[9441]=8'b11111111;
memory[9442]=8'b11111111;
memory[9443]=8'b11111111;
memory[9444]=8'b11111111;
memory[9445]=8'b11111111;
memory[9446]=8'b11111111;
memory[9447]=8'b11111111;
memory[9448]=8'b11111111;
memory[9449]=8'b11111111;
memory[9450]=8'b11111111;
memory[9451]=8'b11111111;
memory[9452]=8'b11111111;
memory[9453]=8'b11111111;
memory[9454]=8'b11111111;
memory[9455]=8'b11111111;
memory[9456]=8'b11111111;
memory[9457]=8'b11111100;
memory[9458]=8'b00000000;
memory[9459]=8'b00000000;
memory[9460]=8'b00111111;
memory[9461]=8'b11111111;
memory[9462]=8'b11111110;
memory[9463]=8'b00111000;
memory[9464]=8'b00011000;
memory[9465]=8'b01000000;
memory[9466]=8'b00111000;
memory[9467]=8'b00111111;
memory[9468]=8'b11111111;
memory[9469]=8'b11001111;
memory[9470]=8'b11111000;
memory[9471]=8'b11111111;
memory[9472]=8'b11111111;
memory[9473]=8'b11111111;
memory[9474]=8'b11111111;
memory[9475]=8'b11111111;
memory[9476]=8'b11111111;
memory[9477]=8'b11111111;
memory[9478]=8'b11111111;
memory[9479]=8'b11111111;
memory[9480]=8'b11111111;
memory[9481]=8'b11111111;
memory[9482]=8'b11111111;
memory[9483]=8'b11111111;
memory[9484]=8'b11111111;
memory[9485]=8'b11111111;
memory[9486]=8'b11111111;
memory[9487]=8'b11111111;
memory[9488]=8'b11111111;
memory[9489]=8'b11111111;
memory[9490]=8'b11111111;
memory[9491]=8'b11111111;
memory[9492]=8'b11111111;
memory[9493]=8'b11111111;
memory[9494]=8'b11111111;
memory[9495]=8'b11111111;
memory[9496]=8'b11111111;
memory[9497]=8'b11111000;
memory[9498]=8'b00000000;
memory[9499]=8'b00000000;
memory[9500]=8'b00011111;
memory[9501]=8'b11111111;
memory[9502]=8'b11111110;
memory[9503]=8'b01110000;
memory[9504]=8'b00010000;
memory[9505]=8'b01100000;
memory[9506]=8'b00111000;
memory[9507]=8'b00001111;
memory[9508]=8'b11111111;
memory[9509]=8'b10001111;
memory[9510]=8'b11111001;
memory[9511]=8'b11111111;
memory[9512]=8'b11111111;
memory[9513]=8'b11111111;
memory[9514]=8'b11111111;
memory[9515]=8'b11111111;
memory[9516]=8'b11111111;
memory[9517]=8'b11111111;
memory[9518]=8'b11111111;
memory[9519]=8'b11111111;
memory[9520]=8'b11111111;
memory[9521]=8'b11111111;
memory[9522]=8'b11111111;
memory[9523]=8'b11111111;
memory[9524]=8'b11111111;
memory[9525]=8'b11111111;
memory[9526]=8'b11111111;
memory[9527]=8'b11111111;
memory[9528]=8'b11111111;
memory[9529]=8'b11111111;
memory[9530]=8'b11111111;
memory[9531]=8'b11111111;
memory[9532]=8'b11111111;
memory[9533]=8'b11111111;
memory[9534]=8'b11111111;
memory[9535]=8'b11111111;
memory[9536]=8'b11111111;
memory[9537]=8'b11110000;
memory[9538]=8'b00000000;
memory[9539]=8'b01111100;
memory[9540]=8'b00011111;
memory[9541]=8'b11111111;
memory[9542]=8'b11111100;
memory[9543]=8'b11110000;
memory[9544]=8'b00000000;
memory[9545]=8'b00110000;
memory[9546]=8'b00000010;
memory[9547]=8'b00000111;
memory[9548]=8'b11111111;
memory[9549]=8'b10011111;
memory[9550]=8'b11111111;
memory[9551]=8'b11111111;
memory[9552]=8'b11111111;
memory[9553]=8'b11111111;
memory[9554]=8'b11111111;
memory[9555]=8'b11111111;
memory[9556]=8'b11111111;
memory[9557]=8'b11111111;
memory[9558]=8'b11111111;
memory[9559]=8'b11111111;
memory[9560]=8'b11111111;
memory[9561]=8'b11111111;
memory[9562]=8'b11111111;
memory[9563]=8'b11111111;
memory[9564]=8'b11111111;
memory[9565]=8'b11111111;
memory[9566]=8'b11111111;
memory[9567]=8'b11111111;
memory[9568]=8'b11111111;
memory[9569]=8'b11111111;
memory[9570]=8'b11111111;
memory[9571]=8'b11111111;
memory[9572]=8'b11111111;
memory[9573]=8'b11111111;
memory[9574]=8'b11111111;
memory[9575]=8'b11111111;
memory[9576]=8'b11111111;
memory[9577]=8'b11100000;
memory[9578]=8'b00000000;
memory[9579]=8'b11101111;
memory[9580]=8'b11111111;
memory[9581]=8'b11111111;
memory[9582]=8'b11111111;
memory[9583]=8'b11100000;
memory[9584]=8'b00000000;
memory[9585]=8'b00110000;
memory[9586]=8'b00000011;
memory[9587]=8'b10000011;
memory[9588]=8'b11111111;
memory[9589]=8'b00011111;
memory[9590]=8'b11111111;
memory[9591]=8'b11111111;
memory[9592]=8'b11111111;
memory[9593]=8'b11111111;
memory[9594]=8'b11111111;
memory[9595]=8'b11111111;
memory[9596]=8'b11111111;
memory[9597]=8'b11111111;
memory[9598]=8'b11111111;
memory[9599]=8'b11111111;
memory[9600]=8'b11111111;
memory[9601]=8'b11111111;
memory[9602]=8'b11111111;
memory[9603]=8'b11111111;
memory[9604]=8'b11111111;
memory[9605]=8'b11111111;
memory[9606]=8'b11111111;
memory[9607]=8'b11111111;
memory[9608]=8'b11111111;
memory[9609]=8'b11111111;
memory[9610]=8'b11111111;
memory[9611]=8'b11111111;
memory[9612]=8'b11111111;
memory[9613]=8'b11111111;
memory[9614]=8'b11111111;
memory[9615]=8'b11111111;
memory[9616]=8'b11111111;
memory[9617]=8'b11000000;
memory[9618]=8'b00000000;
memory[9619]=8'b11111111;
memory[9620]=8'b11111111;
memory[9621]=8'b11111111;
memory[9622]=8'b11111111;
memory[9623]=8'b11100000;
memory[9624]=8'b00100000;
memory[9625]=8'b00111000;
memory[9626]=8'b00011001;
memory[9627]=8'b11110011;
memory[9628]=8'b11111110;
memory[9629]=8'b00111111;
memory[9630]=8'b11111111;
memory[9631]=8'b11111111;
memory[9632]=8'b11111111;
memory[9633]=8'b11111111;
memory[9634]=8'b11111111;
memory[9635]=8'b11111111;
memory[9636]=8'b11111111;
memory[9637]=8'b11111111;
memory[9638]=8'b11111111;
memory[9639]=8'b11111111;
memory[9640]=8'b11111111;
memory[9641]=8'b11111111;
memory[9642]=8'b11111111;
memory[9643]=8'b11111111;
memory[9644]=8'b11111111;
memory[9645]=8'b11111111;
memory[9646]=8'b11111111;
memory[9647]=8'b11111111;
memory[9648]=8'b11111111;
memory[9649]=8'b11111111;
memory[9650]=8'b11111111;
memory[9651]=8'b11111111;
memory[9652]=8'b11111111;
memory[9653]=8'b11111111;
memory[9654]=8'b11111111;
memory[9655]=8'b11111111;
memory[9656]=8'b11111111;
memory[9657]=8'b10000000;
memory[9658]=8'b00000000;
memory[9659]=8'b01111111;
memory[9660]=8'b11111111;
memory[9661]=8'b11111111;
memory[9662]=8'b11111111;
memory[9663]=8'b11100000;
memory[9664]=8'b11000000;
memory[9665]=8'b00111100;
memory[9666]=8'b00111100;
memory[9667]=8'b11111111;
memory[9668]=8'b11111110;
memory[9669]=8'b01111111;
memory[9670]=8'b11111111;
memory[9671]=8'b11111111;
memory[9672]=8'b11111111;
memory[9673]=8'b11111111;
memory[9674]=8'b11111111;
memory[9675]=8'b11111111;
memory[9676]=8'b11111111;
memory[9677]=8'b11111111;
memory[9678]=8'b11111111;
memory[9679]=8'b11111111;
memory[9680]=8'b11111111;
memory[9681]=8'b11111111;
memory[9682]=8'b11111111;
memory[9683]=8'b11111111;
memory[9684]=8'b11111111;
memory[9685]=8'b11111111;
memory[9686]=8'b11111111;
memory[9687]=8'b11111111;
memory[9688]=8'b11111111;
memory[9689]=8'b11111111;
memory[9690]=8'b11111111;
memory[9691]=8'b11111111;
memory[9692]=8'b11111111;
memory[9693]=8'b11111111;
memory[9694]=8'b11111111;
memory[9695]=8'b11111111;
memory[9696]=8'b11111111;
memory[9697]=8'b10000000;
memory[9698]=8'b00000000;
memory[9699]=8'b00001111;
memory[9700]=8'b11111111;
memory[9701]=8'b11111111;
memory[9702]=8'b11111111;
memory[9703]=8'b11110000;
memory[9704]=8'b11000000;
memory[9705]=8'b00011110;
memory[9706]=8'b00111100;
memory[9707]=8'b01111111;
memory[9708]=8'b11111100;
memory[9709]=8'b01111111;
memory[9710]=8'b11111111;
memory[9711]=8'b11111111;
memory[9712]=8'b11111111;
memory[9713]=8'b11111111;
memory[9714]=8'b11111111;
memory[9715]=8'b11111111;
memory[9716]=8'b11111111;
memory[9717]=8'b11111111;
memory[9718]=8'b11111111;
memory[9719]=8'b11111111;
memory[9720]=8'b11111111;
memory[9721]=8'b11111111;
memory[9722]=8'b11111111;
memory[9723]=8'b11111111;
memory[9724]=8'b11111111;
memory[9725]=8'b11111111;
memory[9726]=8'b11111111;
memory[9727]=8'b11111111;
memory[9728]=8'b11111111;
memory[9729]=8'b11111111;
memory[9730]=8'b11111111;
memory[9731]=8'b11111111;
memory[9732]=8'b11111111;
memory[9733]=8'b11111111;
memory[9734]=8'b11111111;
memory[9735]=8'b11111111;
memory[9736]=8'b11111111;
memory[9737]=8'b00000000;
memory[9738]=8'b00000000;
memory[9739]=8'b00000011;
memory[9740]=8'b11111111;
memory[9741]=8'b11111111;
memory[9742]=8'b11111111;
memory[9743]=8'b11110000;
memory[9744]=8'b11100000;
memory[9745]=8'b00011111;
memory[9746]=8'b00111110;
memory[9747]=8'b00111111;
memory[9748]=8'b11111100;
memory[9749]=8'b01111111;
memory[9750]=8'b11111111;
memory[9751]=8'b11111111;
memory[9752]=8'b11111111;
memory[9753]=8'b11111111;
memory[9754]=8'b11111111;
memory[9755]=8'b11111111;
memory[9756]=8'b11111111;
memory[9757]=8'b11111111;
memory[9758]=8'b11111111;
memory[9759]=8'b11111111;
memory[9760]=8'b11111111;
memory[9761]=8'b11111111;
memory[9762]=8'b11111111;
memory[9763]=8'b11111111;
memory[9764]=8'b11111111;
memory[9765]=8'b11111111;
memory[9766]=8'b11111111;
memory[9767]=8'b11111111;
memory[9768]=8'b11111111;
memory[9769]=8'b11111111;
memory[9770]=8'b11111111;
memory[9771]=8'b11111111;
memory[9772]=8'b11111111;
memory[9773]=8'b11111111;
memory[9774]=8'b11111111;
memory[9775]=8'b11111111;
memory[9776]=8'b11111111;
memory[9777]=8'b00000000;
memory[9778]=8'b00000111;
memory[9779]=8'b11100011;
memory[9780]=8'b11111111;
memory[9781]=8'b11111111;
memory[9782]=8'b11111111;
memory[9783]=8'b11111111;
memory[9784]=8'b11110000;
memory[9785]=8'b00111111;
memory[9786]=8'b11111111;
memory[9787]=8'b00011111;
memory[9788]=8'b11111000;
memory[9789]=8'b11111111;
memory[9790]=8'b11111111;
memory[9791]=8'b11111111;
memory[9792]=8'b11111111;
memory[9793]=8'b11111111;
memory[9794]=8'b11111111;
memory[9795]=8'b11111111;
memory[9796]=8'b11111111;
memory[9797]=8'b11111111;
memory[9798]=8'b11111111;
memory[9799]=8'b11111111;
memory[9800]=8'b11111111;
memory[9801]=8'b11111111;
memory[9802]=8'b11111111;
memory[9803]=8'b11111111;
memory[9804]=8'b11111111;
memory[9805]=8'b11111111;
memory[9806]=8'b11111111;
memory[9807]=8'b11111111;
memory[9808]=8'b11111111;
memory[9809]=8'b11111111;
memory[9810]=8'b11111111;
memory[9811]=8'b11111111;
memory[9812]=8'b11111111;
memory[9813]=8'b11111111;
memory[9814]=8'b11111111;
memory[9815]=8'b11111111;
memory[9816]=8'b11111111;
memory[9817]=8'b00000000;
memory[9818]=8'b00011111;
memory[9819]=8'b11111111;
memory[9820]=8'b11111111;
memory[9821]=8'b11111111;
memory[9822]=8'b11111111;
memory[9823]=8'b11111111;
memory[9824]=8'b11111000;
memory[9825]=8'b00011111;
memory[9826]=8'b11111111;
memory[9827]=8'b10001111;
memory[9828]=8'b11110000;
memory[9829]=8'b11111111;
memory[9830]=8'b11111111;
memory[9831]=8'b11111111;
memory[9832]=8'b11111111;
memory[9833]=8'b11111111;
memory[9834]=8'b11111111;
memory[9835]=8'b11111111;
memory[9836]=8'b11111111;
memory[9837]=8'b11111111;
memory[9838]=8'b11111111;
memory[9839]=8'b11111111;
memory[9840]=8'b11111111;
memory[9841]=8'b11111111;
memory[9842]=8'b11111111;
memory[9843]=8'b11111111;
memory[9844]=8'b11111111;
memory[9845]=8'b11111111;
memory[9846]=8'b11111111;
memory[9847]=8'b11111111;
memory[9848]=8'b11111111;
memory[9849]=8'b11111111;
memory[9850]=8'b11111111;
memory[9851]=8'b11111111;
memory[9852]=8'b11111111;
memory[9853]=8'b11111111;
memory[9854]=8'b11111111;
memory[9855]=8'b11111111;
memory[9856]=8'b11111111;
memory[9857]=8'b00000000;
memory[9858]=8'b00111111;
memory[9859]=8'b11111111;
memory[9860]=8'b11111111;
memory[9861]=8'b10101111;
memory[9862]=8'b11111111;
memory[9863]=8'b11111111;
memory[9864]=8'b11111100;
memory[9865]=8'b00111111;
memory[9866]=8'b11111111;
memory[9867]=8'b11001111;
memory[9868]=8'b11110000;
memory[9869]=8'b11111111;
memory[9870]=8'b11111111;
memory[9871]=8'b11111111;
memory[9872]=8'b11111111;
memory[9873]=8'b11111111;
memory[9874]=8'b11111111;
memory[9875]=8'b11111111;
memory[9876]=8'b11111111;
memory[9877]=8'b11111111;
memory[9878]=8'b11111111;
memory[9879]=8'b11111111;
memory[9880]=8'b11111111;
memory[9881]=8'b11111111;
memory[9882]=8'b11111111;
memory[9883]=8'b11111111;
memory[9884]=8'b11111111;
memory[9885]=8'b11111111;
memory[9886]=8'b11111111;
memory[9887]=8'b11111111;
memory[9888]=8'b11111111;
memory[9889]=8'b11111111;
memory[9890]=8'b11111111;
memory[9891]=8'b11111111;
memory[9892]=8'b11111111;
memory[9893]=8'b11111111;
memory[9894]=8'b11111111;
memory[9895]=8'b11111111;
memory[9896]=8'b11111110;
memory[9897]=8'b00000000;
memory[9898]=8'b01111111;
memory[9899]=8'b11111111;
memory[9900]=8'b11111111;
memory[9901]=8'b00000111;
memory[9902]=8'b11111111;
memory[9903]=8'b11111111;
memory[9904]=8'b11111110;
memory[9905]=8'b00111111;
memory[9906]=8'b11111111;
memory[9907]=8'b11000111;
memory[9908]=8'b11100000;
memory[9909]=8'b11111111;
memory[9910]=8'b11111111;
memory[9911]=8'b11111111;
memory[9912]=8'b11111111;
memory[9913]=8'b11111111;
memory[9914]=8'b11111111;
memory[9915]=8'b11111111;
memory[9916]=8'b11111111;
memory[9917]=8'b11111111;
memory[9918]=8'b11111111;
memory[9919]=8'b11111111;
memory[9920]=8'b11111111;
memory[9921]=8'b11111111;
memory[9922]=8'b11111111;
memory[9923]=8'b11111111;
memory[9924]=8'b11111111;
memory[9925]=8'b11111111;
memory[9926]=8'b11111111;
memory[9927]=8'b11111111;
memory[9928]=8'b11111111;
memory[9929]=8'b11111111;
memory[9930]=8'b11111111;
memory[9931]=8'b11111111;
memory[9932]=8'b11111111;
memory[9933]=8'b11111111;
memory[9934]=8'b11111111;
memory[9935]=8'b11111111;
memory[9936]=8'b11111110;
memory[9937]=8'b00000000;
memory[9938]=8'b01111111;
memory[9939]=8'b11111111;
memory[9940]=8'b11111100;
memory[9941]=8'b00000111;
memory[9942]=8'b11111111;
memory[9943]=8'b11111111;
memory[9944]=8'b11111111;
memory[9945]=8'b00111111;
memory[9946]=8'b11111111;
memory[9947]=8'b11100011;
memory[9948]=8'b11100001;
memory[9949]=8'b11111111;
memory[9950]=8'b11111111;
memory[9951]=8'b11111111;
memory[9952]=8'b11111111;
memory[9953]=8'b11111111;
memory[9954]=8'b11111111;
memory[9955]=8'b11111111;
memory[9956]=8'b11111111;
memory[9957]=8'b11111111;
memory[9958]=8'b11111111;
memory[9959]=8'b11111111;
memory[9960]=8'b11111111;
memory[9961]=8'b11111111;
memory[9962]=8'b11111111;
memory[9963]=8'b11111111;
memory[9964]=8'b11111111;
memory[9965]=8'b11111111;
memory[9966]=8'b11111111;
memory[9967]=8'b11111111;
memory[9968]=8'b11111111;
memory[9969]=8'b11111111;
memory[9970]=8'b11111111;
memory[9971]=8'b11111111;
memory[9972]=8'b11111111;
memory[9973]=8'b11111111;
memory[9974]=8'b11111111;
memory[9975]=8'b11111111;
memory[9976]=8'b11111111;
memory[9977]=8'b00000000;
memory[9978]=8'b01111111;
memory[9979]=8'b11111111;
memory[9980]=8'b11111110;
memory[9981]=8'b00001111;
memory[9982]=8'b11111111;
memory[9983]=8'b11111111;
memory[9984]=8'b11111111;
memory[9985]=8'b11111111;
memory[9986]=8'b11111111;
memory[9987]=8'b11100011;
memory[9988]=8'b11000001;
memory[9989]=8'b11111111;
memory[9990]=8'b11111111;
memory[9991]=8'b11111111;
memory[9992]=8'b11111111;
memory[9993]=8'b11111111;
memory[9994]=8'b11111111;
memory[9995]=8'b11111111;
memory[9996]=8'b11111111;
memory[9997]=8'b11111111;
memory[9998]=8'b11111111;
memory[9999]=8'b11111111;
memory[10000]=8'b11111111;
memory[10001]=8'b11111111;
memory[10002]=8'b11111111;
memory[10003]=8'b11111111;
memory[10004]=8'b11111111;
memory[10005]=8'b11111111;
memory[10006]=8'b11111111;
memory[10007]=8'b11111111;
memory[10008]=8'b11111111;
memory[10009]=8'b11111111;
memory[10010]=8'b11111111;
memory[10011]=8'b11111111;
memory[10012]=8'b11111111;
memory[10013]=8'b11111111;
memory[10014]=8'b11111111;
memory[10015]=8'b11111111;
memory[10016]=8'b11111111;
memory[10017]=8'b00000000;
memory[10018]=8'b00111111;
memory[10019]=8'b11111111;
memory[10020]=8'b11111110;
memory[10021]=8'b00001111;
memory[10022]=8'b11111111;
memory[10023]=8'b11111111;
memory[10024]=8'b11111111;
memory[10025]=8'b11111111;
memory[10026]=8'b11111111;
memory[10027]=8'b11110001;
memory[10028]=8'b11000011;
memory[10029]=8'b11111111;
memory[10030]=8'b11111111;
memory[10031]=8'b11111111;
memory[10032]=8'b11111111;
memory[10033]=8'b11111111;
memory[10034]=8'b11111111;
memory[10035]=8'b11111111;
memory[10036]=8'b11111111;
memory[10037]=8'b11111111;
memory[10038]=8'b11111111;
memory[10039]=8'b11111111;
memory[10040]=8'b11111111;
memory[10041]=8'b11111111;
memory[10042]=8'b11111111;
memory[10043]=8'b11111111;
memory[10044]=8'b11111111;
memory[10045]=8'b11111111;
memory[10046]=8'b11111111;
memory[10047]=8'b11111111;
memory[10048]=8'b11111111;
memory[10049]=8'b11111111;
memory[10050]=8'b11111111;
memory[10051]=8'b11111111;
memory[10052]=8'b11111111;
memory[10053]=8'b11111111;
memory[10054]=8'b11111111;
memory[10055]=8'b11111111;
memory[10056]=8'b11111111;
memory[10057]=8'b00000000;
memory[10058]=8'b00011111;
memory[10059]=8'b11111111;
memory[10060]=8'b11111111;
memory[10061]=8'b00001111;
memory[10062]=8'b11111111;
memory[10063]=8'b11111111;
memory[10064]=8'b11111111;
memory[10065]=8'b11111111;
memory[10066]=8'b11111111;
memory[10067]=8'b11110001;
memory[10068]=8'b11000011;
memory[10069]=8'b11111111;
memory[10070]=8'b11111111;
memory[10071]=8'b11111111;
memory[10072]=8'b11111111;
memory[10073]=8'b11111111;
memory[10074]=8'b11111111;
memory[10075]=8'b11111111;
memory[10076]=8'b11111111;
memory[10077]=8'b11111111;
memory[10078]=8'b11111111;
memory[10079]=8'b11111111;
memory[10080]=8'b11111111;
memory[10081]=8'b11111111;
memory[10082]=8'b11111111;
memory[10083]=8'b11111111;
memory[10084]=8'b11111111;
memory[10085]=8'b11111111;
memory[10086]=8'b11111111;
memory[10087]=8'b11111111;
memory[10088]=8'b11111111;
memory[10089]=8'b11111111;
memory[10090]=8'b11111111;
memory[10091]=8'b11111111;
memory[10092]=8'b11111111;
memory[10093]=8'b11111111;
memory[10094]=8'b11111111;
memory[10095]=8'b11111111;
memory[10096]=8'b11111111;
memory[10097]=8'b10000000;
memory[10098]=8'b00001111;
memory[10099]=8'b11111111;
memory[10100]=8'b11111111;
memory[10101]=8'b10001111;
memory[10102]=8'b11111111;
memory[10103]=8'b11111111;
memory[10104]=8'b11111111;
memory[10105]=8'b11111111;
memory[10106]=8'b11111111;
memory[10107]=8'b11110000;
memory[10108]=8'b10000011;
memory[10109]=8'b11111111;
memory[10110]=8'b11111111;
memory[10111]=8'b11111111;
memory[10112]=8'b11111111;
memory[10113]=8'b11111111;
memory[10114]=8'b11111111;
memory[10115]=8'b11111111;
memory[10116]=8'b11111111;
memory[10117]=8'b11111111;
memory[10118]=8'b11111111;
memory[10119]=8'b11111111;
memory[10120]=8'b11111111;
memory[10121]=8'b11111111;
memory[10122]=8'b11111111;
memory[10123]=8'b11111111;
memory[10124]=8'b11111111;
memory[10125]=8'b11111111;
memory[10126]=8'b11111111;
memory[10127]=8'b11111111;
memory[10128]=8'b11111111;
memory[10129]=8'b11111111;
memory[10130]=8'b11111111;
memory[10131]=8'b11111111;
memory[10132]=8'b11111111;
memory[10133]=8'b11111111;
memory[10134]=8'b11111111;
memory[10135]=8'b11111111;
memory[10136]=8'b11111111;
memory[10137]=8'b10000000;
memory[10138]=8'b00001111;
memory[10139]=8'b11111111;
memory[10140]=8'b11111111;
memory[10141]=8'b10011111;
memory[10142]=8'b11111111;
memory[10143]=8'b11111111;
memory[10144]=8'b11111111;
memory[10145]=8'b11111111;
memory[10146]=8'b11111111;
memory[10147]=8'b11111000;
memory[10148]=8'b00000011;
memory[10149]=8'b11111111;
memory[10150]=8'b11111111;
memory[10151]=8'b11111111;
memory[10152]=8'b11111111;
memory[10153]=8'b11111111;
memory[10154]=8'b11111111;
memory[10155]=8'b11111111;
memory[10156]=8'b11111111;
memory[10157]=8'b11111111;
memory[10158]=8'b11111111;
memory[10159]=8'b11111111;
memory[10160]=8'b11111111;
memory[10161]=8'b11111111;
memory[10162]=8'b11111111;
memory[10163]=8'b11111111;
memory[10164]=8'b11111111;
memory[10165]=8'b11111111;
memory[10166]=8'b11111111;
memory[10167]=8'b11111111;
memory[10168]=8'b11111111;
memory[10169]=8'b11111111;
memory[10170]=8'b11111111;
memory[10171]=8'b11111111;
memory[10172]=8'b11111111;
memory[10173]=8'b11111111;
memory[10174]=8'b11111111;
memory[10175]=8'b11111111;
memory[10176]=8'b11111111;
memory[10177]=8'b11000000;
memory[10178]=8'b00000111;
memory[10179]=8'b11111111;
memory[10180]=8'b11111111;
memory[10181]=8'b10011111;
memory[10182]=8'b11111111;
memory[10183]=8'b11111111;
memory[10184]=8'b11111111;
memory[10185]=8'b11111111;
memory[10186]=8'b11111111;
memory[10187]=8'b11111000;
memory[10188]=8'b00000011;
memory[10189]=8'b11111111;
memory[10190]=8'b11111111;
memory[10191]=8'b11111111;
memory[10192]=8'b11111111;
memory[10193]=8'b11111111;
memory[10194]=8'b11111111;
memory[10195]=8'b11111111;
memory[10196]=8'b11111111;
memory[10197]=8'b11111111;
memory[10198]=8'b11111111;
memory[10199]=8'b11111111;
memory[10200]=8'b11111111;
memory[10201]=8'b11111111;
memory[10202]=8'b11111111;
memory[10203]=8'b11111111;
memory[10204]=8'b11111111;
memory[10205]=8'b11111111;
memory[10206]=8'b11111111;
memory[10207]=8'b11111111;
memory[10208]=8'b11111111;
memory[10209]=8'b11111111;
memory[10210]=8'b11111111;
memory[10211]=8'b11111111;
memory[10212]=8'b11111111;
memory[10213]=8'b11111111;
memory[10214]=8'b11111111;
memory[10215]=8'b11111111;
memory[10216]=8'b11111111;
memory[10217]=8'b11100000;
memory[10218]=8'b00000011;
memory[10219]=8'b11111111;
memory[10220]=8'b11111111;
memory[10221]=8'b11111111;
memory[10222]=8'b11111111;
memory[10223]=8'b11111111;
memory[10224]=8'b11111111;
memory[10225]=8'b11111111;
memory[10226]=8'b11111111;
memory[10227]=8'b11110000;
memory[10228]=8'b00100111;
memory[10229]=8'b11111111;
memory[10230]=8'b11111111;
memory[10231]=8'b11111111;
memory[10232]=8'b11111111;
memory[10233]=8'b11111111;
memory[10234]=8'b11111111;
memory[10235]=8'b11111111;
memory[10236]=8'b11111111;
memory[10237]=8'b11111111;
memory[10238]=8'b11111111;
memory[10239]=8'b11111111;
memory[10240]=8'b11111111;
memory[10241]=8'b11111111;
memory[10242]=8'b11111111;
memory[10243]=8'b11111111;
memory[10244]=8'b11111111;
memory[10245]=8'b11111111;
memory[10246]=8'b11111111;
memory[10247]=8'b11111111;
memory[10248]=8'b11111111;
memory[10249]=8'b11111111;
memory[10250]=8'b11111111;
memory[10251]=8'b11111111;
memory[10252]=8'b11111111;
memory[10253]=8'b11111111;
memory[10254]=8'b11111111;
memory[10255]=8'b11111111;
memory[10256]=8'b11111111;
memory[10257]=8'b11100000;
memory[10258]=8'b00000001;
memory[10259]=8'b11111111;
memory[10260]=8'b11111111;
memory[10261]=8'b11111111;
memory[10262]=8'b11111111;
memory[10263]=8'b11111111;
memory[10264]=8'b11111111;
memory[10265]=8'b11111111;
memory[10266]=8'b11111110;
memory[10267]=8'b00000000;
memory[10268]=8'b00000111;
memory[10269]=8'b11111111;
memory[10270]=8'b11111111;
memory[10271]=8'b11111111;
memory[10272]=8'b11111111;
memory[10273]=8'b11111111;
memory[10274]=8'b11111111;
memory[10275]=8'b11111111;
memory[10276]=8'b11111111;
memory[10277]=8'b11111111;
memory[10278]=8'b11111111;
memory[10279]=8'b11111111;
memory[10280]=8'b11111111;
memory[10281]=8'b11111111;
memory[10282]=8'b11111111;
memory[10283]=8'b11111111;
memory[10284]=8'b11111111;
memory[10285]=8'b11111111;
memory[10286]=8'b11111111;
memory[10287]=8'b11111111;
memory[10288]=8'b11111111;
memory[10289]=8'b11111111;
memory[10290]=8'b11111111;
memory[10291]=8'b11111111;
memory[10292]=8'b11111111;
memory[10293]=8'b11111111;
memory[10294]=8'b11111111;
memory[10295]=8'b11111111;
memory[10296]=8'b11111111;
memory[10297]=8'b11110000;
memory[10298]=8'b00000000;
memory[10299]=8'b11111111;
memory[10300]=8'b11111111;
memory[10301]=8'b11111111;
memory[10302]=8'b11111111;
memory[10303]=8'b11111111;
memory[10304]=8'b11111111;
memory[10305]=8'b11111111;
memory[10306]=8'b11110000;
memory[10307]=8'b00000000;
memory[10308]=8'b00000000;
memory[10309]=8'b11111111;
memory[10310]=8'b11111111;
memory[10311]=8'b11111111;
memory[10312]=8'b11111111;
memory[10313]=8'b11111111;
memory[10314]=8'b11111111;
memory[10315]=8'b11111111;
memory[10316]=8'b11111111;
memory[10317]=8'b11111111;
memory[10318]=8'b11111111;
memory[10319]=8'b11111111;
memory[10320]=8'b11111111;
memory[10321]=8'b11111111;
memory[10322]=8'b11111111;
memory[10323]=8'b11111111;
memory[10324]=8'b11111111;
memory[10325]=8'b11111111;
memory[10326]=8'b11111111;
memory[10327]=8'b11111111;
memory[10328]=8'b11111111;
memory[10329]=8'b11111111;
memory[10330]=8'b11111111;
memory[10331]=8'b11111111;
memory[10332]=8'b11111111;
memory[10333]=8'b11111111;
memory[10334]=8'b11111111;
memory[10335]=8'b11111111;
memory[10336]=8'b11111111;
memory[10337]=8'b11111000;
memory[10338]=8'b00000000;
memory[10339]=8'b01111111;
memory[10340]=8'b11111111;
memory[10341]=8'b11111111;
memory[10342]=8'b11111111;
memory[10343]=8'b11111111;
memory[10344]=8'b11111111;
memory[10345]=8'b11111111;
memory[10346]=8'b10000000;
memory[10347]=8'b00000000;
memory[10348]=8'b00000000;
memory[10349]=8'b00011111;
memory[10350]=8'b11111111;
memory[10351]=8'b11111111;
memory[10352]=8'b11111111;
memory[10353]=8'b11111111;
memory[10354]=8'b11111111;
memory[10355]=8'b11111111;
memory[10356]=8'b11111111;
memory[10357]=8'b11111111;
memory[10358]=8'b11111111;
memory[10359]=8'b11111111;
memory[10360]=8'b11111111;
memory[10361]=8'b11111111;
memory[10362]=8'b11111111;
memory[10363]=8'b11111111;
memory[10364]=8'b11111111;
memory[10365]=8'b11111111;
memory[10366]=8'b11111111;
memory[10367]=8'b11111111;
memory[10368]=8'b00000000;
memory[10369]=8'b00000000;
memory[10370]=8'b00000000;
memory[10371]=8'b00000000;
memory[10372]=8'b00000000;
memory[10373]=8'b00000000;
memory[10374]=8'b00000000;
memory[10375]=8'b00000000;
memory[10376]=8'b00000111;
memory[10377]=8'b11111100;
memory[10378]=8'b00000000;
memory[10379]=8'b00111111;
memory[10380]=8'b11111111;
memory[10381]=8'b11000000;
memory[10382]=8'b00000000;
memory[10383]=8'b00111111;
memory[10384]=8'b11111111;
memory[10385]=8'b11111110;
memory[10386]=8'b00000000;
memory[10387]=8'b00000000;
memory[10388]=8'b00000000;
memory[10389]=8'b00000111;
memory[10390]=8'b11111111;
memory[10391]=8'b11111111;
memory[10392]=8'b11111111;
memory[10393]=8'b11111111;
memory[10394]=8'b11111111;
memory[10395]=8'b11111111;
memory[10396]=8'b11111111;
memory[10397]=8'b11111111;
memory[10398]=8'b11111111;
memory[10399]=8'b11111111;
memory[10400]=8'b11111111;
memory[10401]=8'b11111111;
memory[10402]=8'b11111111;
memory[10403]=8'b11111111;
memory[10404]=8'b11111111;
memory[10405]=8'b11111111;
memory[10406]=8'b11111111;
memory[10407]=8'b11111111;
memory[10408]=8'b11110000;
memory[10409]=8'b00000000;
memory[10410]=8'b01111111;
memory[10411]=8'b11111110;
memory[10412]=8'b00000000;
memory[10413]=8'b01111111;
memory[10414]=8'b11111100;
memory[10415]=8'b00000111;
memory[10416]=8'b11111111;
memory[10417]=8'b11111110;
memory[10418]=8'b00000000;
memory[10419]=8'b00011111;
memory[10420]=8'b11111111;
memory[10421]=8'b11111111;
memory[10422]=8'b11111111;
memory[10423]=8'b11111111;
memory[10424]=8'b11111111;
memory[10425]=8'b11110000;
memory[10426]=8'b00000000;
memory[10427]=8'b00000000;
memory[10428]=8'b00000000;
memory[10429]=8'b00000001;
memory[10430]=8'b11111111;
memory[10431]=8'b11111111;
memory[10432]=8'b11111111;
memory[10433]=8'b11111111;
memory[10434]=8'b11111111;
memory[10435]=8'b11111111;
memory[10436]=8'b11111111;
memory[10437]=8'b11111111;
memory[10438]=8'b11111111;
memory[10439]=8'b11111111;
memory[10440]=8'b11111111;
memory[10441]=8'b11111111;
memory[10442]=8'b11111111;
memory[10443]=8'b11111111;
memory[10444]=8'b11111111;
memory[10445]=8'b11111111;
memory[10446]=8'b11111111;
memory[10447]=8'b11111111;
memory[10448]=8'b11111111;
memory[10449]=8'b11111111;
memory[10450]=8'b11111111;
memory[10451]=8'b11111111;
memory[10452]=8'b11111111;
memory[10453]=8'b11111111;
memory[10454]=8'b11111111;
memory[10455]=8'b11111111;
memory[10456]=8'b11111111;
memory[10457]=8'b11111111;
memory[10458]=8'b00000000;
memory[10459]=8'b00001111;
memory[10460]=8'b11111111;
memory[10461]=8'b11111111;
memory[10462]=8'b11111111;
memory[10463]=8'b11111111;
memory[10464]=8'b11111111;
memory[10465]=8'b00000000;
memory[10466]=8'b00000000;
memory[10467]=8'b00000000;
memory[10468]=8'b00000000;
memory[10469]=8'b00000000;
memory[10470]=8'b01111111;
memory[10471]=8'b11111111;
memory[10472]=8'b11111111;
memory[10473]=8'b11111111;
memory[10474]=8'b11111111;
memory[10475]=8'b11111111;
memory[10476]=8'b11111111;
memory[10477]=8'b11111111;
memory[10478]=8'b11111111;
memory[10479]=8'b11111111;
memory[10480]=8'b11111111;
memory[10481]=8'b11111111;
memory[10482]=8'b11111111;
memory[10483]=8'b11111111;
memory[10484]=8'b11111111;
memory[10485]=8'b11111111;
memory[10486]=8'b11111111;
memory[10487]=8'b11111111;
memory[10488]=8'b11111111;
memory[10489]=8'b11111111;
memory[10490]=8'b11111111;
memory[10491]=8'b11111111;
memory[10492]=8'b11111111;
memory[10493]=8'b11111111;
memory[10494]=8'b11111111;
memory[10495]=8'b11111111;
memory[10496]=8'b11111111;
memory[10497]=8'b11111111;
memory[10498]=8'b11000000;
memory[10499]=8'b00000111;
memory[10500]=8'b11111111;
memory[10501]=8'b11111111;
memory[10502]=8'b11111111;
memory[10503]=8'b11111111;
memory[10504]=8'b11110000;
memory[10505]=8'b00000000;
memory[10506]=8'b00000000;
memory[10507]=8'b00000000;
memory[10508]=8'b00000000;
memory[10509]=8'b00000000;
memory[10510]=8'b00011111;
memory[10511]=8'b11111111;
memory[10512]=8'b11111111;
memory[10513]=8'b11111111;
memory[10514]=8'b11111111;
memory[10515]=8'b11111111;
memory[10516]=8'b11111111;
memory[10517]=8'b11111111;
memory[10518]=8'b11111111;
memory[10519]=8'b11111111;
memory[10520]=8'b11111111;
memory[10521]=8'b11111111;
memory[10522]=8'b11111111;
memory[10523]=8'b11111111;
memory[10524]=8'b11111111;
memory[10525]=8'b11111111;
memory[10526]=8'b11111111;
memory[10527]=8'b11111111;
memory[10528]=8'b11111111;
memory[10529]=8'b11111111;
memory[10530]=8'b11111111;
memory[10531]=8'b11111111;
memory[10532]=8'b11111111;
memory[10533]=8'b11111111;
memory[10534]=8'b11111111;
memory[10535]=8'b11111111;
memory[10536]=8'b11111111;
memory[10537]=8'b11111111;
memory[10538]=8'b11100000;
memory[10539]=8'b00000011;
memory[10540]=8'b11111111;
memory[10541]=8'b11111111;
memory[10542]=8'b11111111;
memory[10543]=8'b11111111;
memory[10544]=8'b10000000;
memory[10545]=8'b00000000;
memory[10546]=8'b00000000;
memory[10547]=8'b00000000;
memory[10548]=8'b00000000;
memory[10549]=8'b00000000;
memory[10550]=8'b00000001;
memory[10551]=8'b11111111;
memory[10552]=8'b11111111;
memory[10553]=8'b11111111;
memory[10554]=8'b11111111;
memory[10555]=8'b11111111;
memory[10556]=8'b11111111;
memory[10557]=8'b11111111;
memory[10558]=8'b11111111;
memory[10559]=8'b11111111;
memory[10560]=8'b11111111;
memory[10561]=8'b11111111;
memory[10562]=8'b11111111;
memory[10563]=8'b11111111;
memory[10564]=8'b11111111;
memory[10565]=8'b11111111;
memory[10566]=8'b11111111;
memory[10567]=8'b11111111;
memory[10568]=8'b11111111;
memory[10569]=8'b11111111;
memory[10570]=8'b11111111;
memory[10571]=8'b11111111;
memory[10572]=8'b11111111;
memory[10573]=8'b11111111;
memory[10574]=8'b11111111;
memory[10575]=8'b11111111;
memory[10576]=8'b11111111;
memory[10577]=8'b11111111;
memory[10578]=8'b11110000;
memory[10579]=8'b00000001;
memory[10580]=8'b11111111;
memory[10581]=8'b11111111;
memory[10582]=8'b11111111;
memory[10583]=8'b11111111;
memory[10584]=8'b10001111;
memory[10585]=8'b10000000;
memory[10586]=8'b00000000;
memory[10587]=8'b00000000;
memory[10588]=8'b00111000;
memory[10589]=8'b00000000;
memory[10590]=8'b00000000;
memory[10591]=8'b01111111;
memory[10592]=8'b11111111;
memory[10593]=8'b11111111;
memory[10594]=8'b11111111;
memory[10595]=8'b11111111;
memory[10596]=8'b11111111;
memory[10597]=8'b11111111;
memory[10598]=8'b11111111;
memory[10599]=8'b11111111;
memory[10600]=8'b11111111;
memory[10601]=8'b11111111;
memory[10602]=8'b11111111;
memory[10603]=8'b11111111;
memory[10604]=8'b11111111;
memory[10605]=8'b11111111;
memory[10606]=8'b11111111;
memory[10607]=8'b11111111;
memory[10608]=8'b11111111;
memory[10609]=8'b11111111;
memory[10610]=8'b11111111;
memory[10611]=8'b11111111;
memory[10612]=8'b11111111;
memory[10613]=8'b11111111;
memory[10614]=8'b11111111;
memory[10615]=8'b11111111;
memory[10616]=8'b11111111;
memory[10617]=8'b11111111;
memory[10618]=8'b11111000;
memory[10619]=8'b00000000;
memory[10620]=8'b11111111;
memory[10621]=8'b11111111;
memory[10622]=8'b11111111;
memory[10623]=8'b11111111;
memory[10624]=8'b11111111;
memory[10625]=8'b11111100;
memory[10626]=8'b00000000;
memory[10627]=8'b11111111;
memory[10628]=8'b11111111;
memory[10629]=8'b11111111;
memory[10630]=8'b11111111;
memory[10631]=8'b11111111;
memory[10632]=8'b11111111;
memory[10633]=8'b11111111;
memory[10634]=8'b11111111;
memory[10635]=8'b11111111;
memory[10636]=8'b11111111;
memory[10637]=8'b11111111;
memory[10638]=8'b11111111;
memory[10639]=8'b11111111;
memory[10640]=8'b11111111;
memory[10641]=8'b11111111;
memory[10642]=8'b11111111;
memory[10643]=8'b11111111;
memory[10644]=8'b11111111;
memory[10645]=8'b11111111;
memory[10646]=8'b11111111;
memory[10647]=8'b11111111;
memory[10648]=8'b11111111;
memory[10649]=8'b11111111;
memory[10650]=8'b11111111;
memory[10651]=8'b11111111;
memory[10652]=8'b11111111;
memory[10653]=8'b11111111;
memory[10654]=8'b11111111;
memory[10655]=8'b11111111;
memory[10656]=8'b11111111;
memory[10657]=8'b11111111;
memory[10658]=8'b11111100;
memory[10659]=8'b00000000;
memory[10660]=8'b01111111;
memory[10661]=8'b11111111;
memory[10662]=8'b11111111;
memory[10663]=8'b11111111;
memory[10664]=8'b11111111;
memory[10665]=8'b11111111;
memory[10666]=8'b11111111;
memory[10667]=8'b11111111;
memory[10668]=8'b11111111;
memory[10669]=8'b11111111;
memory[10670]=8'b11111111;
memory[10671]=8'b11111111;
memory[10672]=8'b11111111;
memory[10673]=8'b11111111;
memory[10674]=8'b11111111;
memory[10675]=8'b11111111;
memory[10676]=8'b11111111;
memory[10677]=8'b11111111;
memory[10678]=8'b11111111;
memory[10679]=8'b11111111;
memory[10680]=8'b11111111;
memory[10681]=8'b11111111;
memory[10682]=8'b11111111;
memory[10683]=8'b11111111;
memory[10684]=8'b11111111;
memory[10685]=8'b11111111;
memory[10686]=8'b11111111;
memory[10687]=8'b11111111;
memory[10688]=8'b11111111;
memory[10689]=8'b11111111;
memory[10690]=8'b11111111;
memory[10691]=8'b11111111;
memory[10692]=8'b11111111;
memory[10693]=8'b11111111;
memory[10694]=8'b11111111;
memory[10695]=8'b11111111;
memory[10696]=8'b11111111;
memory[10697]=8'b11111111;
memory[10698]=8'b11111110;
memory[10699]=8'b00000000;
memory[10700]=8'b00111111;
memory[10701]=8'b11111111;
memory[10702]=8'b11111111;
memory[10703]=8'b11111111;
memory[10704]=8'b11111111;
memory[10705]=8'b11111111;
memory[10706]=8'b11111111;
memory[10707]=8'b11111111;
memory[10708]=8'b11111111;
memory[10709]=8'b11111111;
memory[10710]=8'b11111111;
memory[10711]=8'b11111111;
memory[10712]=8'b11111111;
memory[10713]=8'b11111111;
memory[10714]=8'b11111111;
memory[10715]=8'b11111111;
memory[10716]=8'b11111111;
memory[10717]=8'b11111111;
memory[10718]=8'b11111111;
memory[10719]=8'b11111111;
memory[10720]=8'b11111111;
memory[10721]=8'b11111111;
memory[10722]=8'b11111111;
memory[10723]=8'b11111111;
memory[10724]=8'b11111111;
memory[10725]=8'b11111111;
memory[10726]=8'b11111111;
memory[10727]=8'b11111111;
memory[10728]=8'b11111111;
memory[10729]=8'b11111111;
memory[10730]=8'b11111111;
memory[10731]=8'b11111111;
memory[10732]=8'b11111111;
memory[10733]=8'b11111111;
memory[10734]=8'b10000000;
memory[10735]=8'b00111111;
memory[10736]=8'b11111111;
memory[10737]=8'b11111111;
memory[10738]=8'b11111111;
memory[10739]=8'b10000000;
memory[10740]=8'b00111111;
memory[10741]=8'b11111111;
memory[10742]=8'b11111111;
memory[10743]=8'b11111111;
memory[10744]=8'b11111111;
memory[10745]=8'b11111111;
memory[10746]=8'b11111111;
memory[10747]=8'b11111111;
memory[10748]=8'b11100000;
memory[10749]=8'b00000000;
memory[10750]=8'b00000000;
memory[10751]=8'b00000000;
memory[10752]=8'b01111111;
memory[10753]=8'b11111111;
memory[10754]=8'b11111111;
memory[10755]=8'b11111111;
memory[10756]=8'b11111111;
memory[10757]=8'b11111111;
memory[10758]=8'b11111111;
memory[10759]=8'b11111111;
memory[10760]=8'b11111111;
memory[10761]=8'b11111111;
memory[10762]=8'b11111111;
memory[10763]=8'b11111111;
memory[10764]=8'b11111111;
memory[10765]=8'b11111111;
memory[10766]=8'b11111111;
memory[10767]=8'b11111111;
memory[10768]=8'b11111111;
memory[10769]=8'b11111111;
memory[10770]=8'b11111111;
memory[10771]=8'b11111111;
memory[10772]=8'b11111111;
memory[10773]=8'b00000000;
memory[10774]=8'b00000000;
memory[10775]=8'b00000000;
memory[10776]=8'b01111111;
memory[10777]=8'b11111111;
memory[10778]=8'b11111111;
memory[10779]=8'b10000000;
memory[10780]=8'b00011111;
memory[10781]=8'b11111111;
memory[10782]=8'b11111111;
memory[10783]=8'b11111111;
memory[10784]=8'b11111111;
memory[10785]=8'b11111111;
memory[10786]=8'b11111111;
memory[10787]=8'b11111111;
memory[10788]=8'b11111111;
memory[10789]=8'b11000000;
memory[10790]=8'b00000111;
memory[10791]=8'b11111111;
memory[10792]=8'b11111111;
memory[10793]=8'b11111111;
memory[10794]=8'b11111111;
memory[10795]=8'b11111111;
memory[10796]=8'b11111111;
memory[10797]=8'b11111111;
memory[10798]=8'b11111111;
memory[10799]=8'b11111111;
memory[10800]=8'b11111111;
memory[10801]=8'b11111111;
memory[10802]=8'b11111111;
memory[10803]=8'b11111111;
memory[10804]=8'b11111111;
memory[10805]=8'b11111111;
memory[10806]=8'b11111111;
memory[10807]=8'b11111111;
memory[10808]=8'b11111111;
memory[10809]=8'b11111111;
memory[10810]=8'b11111111;
memory[10811]=8'b11111111;
memory[10812]=8'b11111111;
memory[10813]=8'b11111111;
memory[10814]=8'b11110000;
memory[10815]=8'b00000000;
memory[10816]=8'b00001111;
memory[10817]=8'b11111111;
memory[10818]=8'b11111111;
memory[10819]=8'b11000000;
memory[10820]=8'b00001111;
memory[10821]=8'b11111111;
memory[10822]=8'b11111111;
memory[10823]=8'b11111111;
memory[10824]=8'b11111111;
memory[10825]=8'b11111111;
memory[10826]=8'b11101111;
memory[10827]=8'b11111100;
memory[10828]=8'b00011000;
memory[10829]=8'b00000000;
memory[10830]=8'b00000011;
memory[10831]=8'b11111111;
memory[10832]=8'b11111111;
memory[10833]=8'b11111111;
memory[10834]=8'b11111111;
memory[10835]=8'b11111111;
memory[10836]=8'b11111111;
memory[10837]=8'b11111111;
memory[10838]=8'b11111111;
memory[10839]=8'b11111111;
memory[10840]=8'b11111111;
memory[10841]=8'b11111111;
memory[10842]=8'b11111111;
memory[10843]=8'b11111111;
memory[10844]=8'b11111111;
memory[10845]=8'b11111111;
memory[10846]=8'b11111111;
memory[10847]=8'b11111111;
memory[10848]=8'b11111111;
memory[10849]=8'b11111111;
memory[10850]=8'b11111111;
memory[10851]=8'b11111000;
memory[10852]=8'b00111111;
memory[10853]=8'b11111111;
memory[10854]=8'b11111111;
memory[10855]=8'b10000000;
memory[10856]=8'b00000001;
memory[10857]=8'b11111111;
memory[10858]=8'b11111111;
memory[10859]=8'b11100000;
memory[10860]=8'b00000111;
memory[10861]=8'b11111111;
memory[10862]=8'b11111111;
memory[10863]=8'b11111111;
memory[10864]=8'b11111111;
memory[10865]=8'b11111111;
memory[10866]=8'b11111111;
memory[10867]=8'b11111111;
memory[10868]=8'b11100000;
memory[10869]=8'b00000000;
memory[10870]=8'b00000011;
memory[10871]=8'b11111111;
memory[10872]=8'b11111111;
memory[10873]=8'b11111111;
memory[10874]=8'b11111111;
memory[10875]=8'b11111111;
memory[10876]=8'b11111111;
memory[10877]=8'b11111111;
memory[10878]=8'b11111111;
memory[10879]=8'b11111111;
memory[10880]=8'b11111111;
memory[10881]=8'b11111111;
memory[10882]=8'b11111111;
memory[10883]=8'b11111111;
memory[10884]=8'b11111111;
memory[10885]=8'b11111111;
memory[10886]=8'b11111111;
memory[10887]=8'b11111111;
memory[10888]=8'b11111111;
memory[10889]=8'b11111111;
memory[10890]=8'b11111111;
memory[10891]=8'b11000001;
memory[10892]=8'b11111111;
memory[10893]=8'b11111111;
memory[10894]=8'b11111100;
memory[10895]=8'b00000000;
memory[10896]=8'b00000000;
memory[10897]=8'b01111111;
memory[10898]=8'b11111111;
memory[10899]=8'b11110000;
memory[10900]=8'b00000111;
memory[10901]=8'b11111111;
memory[10902]=8'b11111111;
memory[10903]=8'b11111111;
memory[10904]=8'b11111111;
memory[10905]=8'b11111111;
memory[10906]=8'b11111111;
memory[10907]=8'b11111111;
memory[10908]=8'b11100000;
memory[10909]=8'b00000000;
memory[10910]=8'b00001111;
memory[10911]=8'b11111111;
memory[10912]=8'b11111111;
memory[10913]=8'b11111111;
memory[10914]=8'b11111111;
memory[10915]=8'b11111111;
memory[10916]=8'b11111111;
memory[10917]=8'b11111111;
memory[10918]=8'b11111111;
memory[10919]=8'b11111111;
memory[10920]=8'b11111111;
memory[10921]=8'b11111111;
memory[10922]=8'b11111111;
memory[10923]=8'b11111111;
memory[10924]=8'b11111111;
memory[10925]=8'b11111111;
memory[10926]=8'b11111111;
memory[10927]=8'b11111111;
memory[10928]=8'b11111111;
memory[10929]=8'b11111111;
memory[10930]=8'b11111110;
memory[10931]=8'b00001111;
memory[10932]=8'b11111111;
memory[10933]=8'b11111111;
memory[10934]=8'b11111111;
memory[10935]=8'b11100000;
memory[10936]=8'b00000000;
memory[10937]=8'b00011111;
memory[10938]=8'b11111111;
memory[10939]=8'b11111000;
memory[10940]=8'b00000011;
memory[10941]=8'b11111111;
memory[10942]=8'b11111111;
memory[10943]=8'b11100001;
memory[10944]=8'b11111111;
memory[10945]=8'b11111111;
memory[10946]=8'b11100000;
memory[10947]=8'b00000000;
memory[10948]=8'b00000000;
memory[10949]=8'b00000000;
memory[10950]=8'b00000000;
memory[10951]=8'b00000000;
memory[10952]=8'b00011111;
memory[10953]=8'b11111111;
memory[10954]=8'b11111111;
memory[10955]=8'b11111111;
memory[10956]=8'b11111111;
memory[10957]=8'b11111111;
memory[10958]=8'b11111111;
memory[10959]=8'b11111111;
memory[10960]=8'b11111111;
memory[10961]=8'b11111111;
memory[10962]=8'b11111111;
memory[10963]=8'b11111111;
memory[10964]=8'b11111111;
memory[10965]=8'b11111111;
memory[10966]=8'b11111111;
memory[10967]=8'b11111111;
memory[10968]=8'b11111111;
memory[10969]=8'b11111111;
memory[10970]=8'b11110000;
memory[10971]=8'b00111111;
memory[10972]=8'b11111111;
memory[10973]=8'b11101111;
memory[10974]=8'b11111111;
memory[10975]=8'b11111000;
memory[10976]=8'b00000000;
memory[10977]=8'b00001111;
memory[10978]=8'b11111111;
memory[10979]=8'b11111000;
memory[10980]=8'b00000001;
memory[10981]=8'b11111111;
memory[10982]=8'b11111100;
memory[10983]=8'b00000000;
memory[10984]=8'b00011111;
memory[10985]=8'b11111111;
memory[10986]=8'b11111111;
memory[10987]=8'b11111110;
memory[10988]=8'b00000000;
memory[10989]=8'b00000000;
memory[10990]=8'b00001111;
memory[10991]=8'b11111111;
memory[10992]=8'b11111111;
memory[10993]=8'b11111111;
memory[10994]=8'b11111111;
memory[10995]=8'b11111111;
memory[10996]=8'b11111111;
memory[10997]=8'b11111111;
memory[10998]=8'b11111111;
memory[10999]=8'b11111111;
memory[11000]=8'b11111111;
memory[11001]=8'b11111111;
memory[11002]=8'b11111111;
memory[11003]=8'b11111111;
memory[11004]=8'b11111111;
memory[11005]=8'b11111111;
memory[11006]=8'b11111111;
memory[11007]=8'b11111111;
memory[11008]=8'b11111111;
memory[11009]=8'b11111111;
memory[11010]=8'b11100011;
memory[11011]=8'b11111111;
memory[11012]=8'b11111111;
memory[11013]=8'b10011111;
memory[11014]=8'b11111111;
memory[11015]=8'b11111100;
memory[11016]=8'b00000000;
memory[11017]=8'b00000111;
memory[11018]=8'b11111111;
memory[11019]=8'b11111100;
memory[11020]=8'b00000001;
memory[11021]=8'b11111111;
memory[11022]=8'b11111000;
memory[11023]=8'b00000000;
memory[11024]=8'b00000111;
memory[11025]=8'b11111111;
memory[11026]=8'b11111111;
memory[11027]=8'b11111111;
memory[11028]=8'b11100000;
memory[11029]=8'b00000000;
memory[11030]=8'b00000111;
memory[11031]=8'b11111111;
memory[11032]=8'b11111111;
memory[11033]=8'b11111111;
memory[11034]=8'b11111111;
memory[11035]=8'b11111111;
memory[11036]=8'b11111111;
memory[11037]=8'b11111111;
memory[11038]=8'b11111111;
memory[11039]=8'b11111111;
memory[11040]=8'b11111111;
memory[11041]=8'b11111111;
memory[11042]=8'b11111111;
memory[11043]=8'b11111111;
memory[11044]=8'b11111111;
memory[11045]=8'b11111111;
memory[11046]=8'b11111111;
memory[11047]=8'b11111111;
memory[11048]=8'b11111111;
memory[11049]=8'b11111111;
memory[11050]=8'b10011111;
memory[11051]=8'b11111111;
memory[11052]=8'b11111111;
memory[11053]=8'b00011111;
memory[11054]=8'b10111111;
memory[11055]=8'b11111100;
memory[11056]=8'b00000000;
memory[11057]=8'b00000011;
memory[11058]=8'b11111111;
memory[11059]=8'b11111110;
memory[11060]=8'b00000000;
memory[11061]=8'b11111111;
memory[11062]=8'b11111000;
memory[11063]=8'b01111000;
memory[11064]=8'b00000011;
memory[11065]=8'b11111111;
memory[11066]=8'b11100000;
memory[11067]=8'b00011111;
memory[11068]=8'b11000000;
memory[11069]=8'b00000000;
memory[11070]=8'b11111111;
memory[11071]=8'b11111111;
memory[11072]=8'b11111111;
memory[11073]=8'b11111111;
memory[11074]=8'b11111111;
memory[11075]=8'b11111111;
memory[11076]=8'b11111111;
memory[11077]=8'b11111111;
memory[11078]=8'b11111111;
memory[11079]=8'b11111111;
memory[11080]=8'b11111111;
memory[11081]=8'b11111111;
memory[11082]=8'b11111111;
memory[11083]=8'b11111111;
memory[11084]=8'b11111111;
memory[11085]=8'b11111111;
memory[11086]=8'b11111111;
memory[11087]=8'b11111111;
memory[11088]=8'b11111111;
memory[11089]=8'b11111110;
memory[11090]=8'b01111111;
memory[11091]=8'b11111111;
memory[11092]=8'b11111111;
memory[11093]=8'b00011110;
memory[11094]=8'b00111111;
memory[11095]=8'b11111000;
memory[11096]=8'b00000000;
memory[11097]=8'b00000001;
memory[11098]=8'b11111111;
memory[11099]=8'b11111110;
memory[11100]=8'b00000000;
memory[11101]=8'b11111111;
memory[11102]=8'b11111111;
memory[11103]=8'b11111100;
memory[11104]=8'b00000001;
memory[11105]=8'b11111111;
memory[11106]=8'b11100000;
memory[11107]=8'b01111111;
memory[11108]=8'b11111000;
memory[11109]=8'b00000111;
memory[11110]=8'b11111111;
memory[11111]=8'b11111111;
memory[11112]=8'b11111111;
memory[11113]=8'b11111111;
memory[11114]=8'b11111111;
memory[11115]=8'b11111111;
memory[11116]=8'b11111111;
memory[11117]=8'b11111111;
memory[11118]=8'b11111111;
memory[11119]=8'b11111111;
memory[11120]=8'b11111111;
memory[11121]=8'b11111111;
memory[11122]=8'b11111111;
memory[11123]=8'b11111111;
memory[11124]=8'b11111111;
memory[11125]=8'b11111111;
memory[11126]=8'b11111111;
memory[11127]=8'b11111111;
memory[11128]=8'b11111111;
memory[11129]=8'b11111111;
memory[11130]=8'b11111111;
memory[11131]=8'b11101111;
memory[11132]=8'b11111111;
memory[11133]=8'b00000000;
memory[11134]=8'b01111111;
memory[11135]=8'b11100000;
memory[11136]=8'b00000000;
memory[11137]=8'b00000000;
memory[11138]=8'b11111111;
memory[11139]=8'b11111110;
memory[11140]=8'b00000000;
memory[11141]=8'b11111111;
memory[11142]=8'b11111111;
memory[11143]=8'b11110000;
memory[11144]=8'b00000000;
memory[11145]=8'b11111111;
memory[11146]=8'b11111111;
memory[11147]=8'b11111111;
memory[11148]=8'b11111100;
memory[11149]=8'b00000011;
memory[11150]=8'b11111111;
memory[11151]=8'b11111111;
memory[11152]=8'b11111111;
memory[11153]=8'b11111111;
memory[11154]=8'b11111111;
memory[11155]=8'b11111111;
memory[11156]=8'b11111111;
memory[11157]=8'b11111111;
memory[11158]=8'b11111111;
memory[11159]=8'b11111111;
memory[11160]=8'b11111111;
memory[11161]=8'b11111111;
memory[11162]=8'b11111111;
memory[11163]=8'b11111111;
memory[11164]=8'b11111111;
memory[11165]=8'b11111111;
memory[11166]=8'b11111111;
memory[11167]=8'b11111111;
memory[11168]=8'b11111111;
memory[11169]=8'b11111111;
memory[11170]=8'b11111111;
memory[11171]=8'b11011111;
memory[11172]=8'b11111111;
memory[11173]=8'b00000000;
memory[11174]=8'b01111111;
memory[11175]=8'b11111110;
memory[11176]=8'b00000000;
memory[11177]=8'b00000000;
memory[11178]=8'b01111111;
memory[11179]=8'b11111110;
memory[11180]=8'b00000000;
memory[11181]=8'b01111111;
memory[11182]=8'b11111111;
memory[11183]=8'b11000000;
memory[11184]=8'b00000000;
memory[11185]=8'b01111111;
memory[11186]=8'b11111111;
memory[11187]=8'b11100000;
memory[11188]=8'b00000000;
memory[11189]=8'b00000000;
memory[11190]=8'b00000000;
memory[11191]=8'b01111111;
memory[11192]=8'b11111111;
memory[11193]=8'b11111111;
memory[11194]=8'b11111111;
memory[11195]=8'b11111111;
memory[11196]=8'b11111111;
memory[11197]=8'b11111111;
memory[11198]=8'b11111111;
memory[11199]=8'b11111111;
memory[11200]=8'b11111111;
memory[11201]=8'b11111111;
memory[11202]=8'b11111111;
memory[11203]=8'b11111111;
memory[11204]=8'b11111111;
memory[11205]=8'b11111111;
memory[11206]=8'b11111111;
memory[11207]=8'b11111111;
memory[11208]=8'b11111111;
memory[11209]=8'b11111111;
memory[11210]=8'b11111111;
memory[11211]=8'b10011111;
memory[11212]=8'b11110010;
memory[11213]=8'b00000000;
memory[11214]=8'b00011111;
memory[11215]=8'b11111111;
memory[11216]=8'b00000000;
memory[11217]=8'b00000000;
memory[11218]=8'b01111111;
memory[11219]=8'b11111111;
memory[11220]=8'b00000000;
memory[11221]=8'b01111111;
memory[11222]=8'b11111111;
memory[11223]=8'b00000000;
memory[11224]=8'b00000000;
memory[11225]=8'b01111111;
memory[11226]=8'b11111111;
memory[11227]=8'b11110000;
memory[11228]=8'b00000011;
memory[11229]=8'b11111111;
memory[11230]=8'b11111111;
memory[11231]=8'b11111111;
memory[11232]=8'b11111111;
memory[11233]=8'b11111111;
memory[11234]=8'b11111111;
memory[11235]=8'b11111111;
memory[11236]=8'b11111111;
memory[11237]=8'b11111111;
memory[11238]=8'b11111111;
memory[11239]=8'b11111111;
memory[11240]=8'b11111111;
memory[11241]=8'b11111111;
memory[11242]=8'b11111111;
memory[11243]=8'b11111111;
memory[11244]=8'b11111111;
memory[11245]=8'b11111111;
memory[11246]=8'b11111111;
memory[11247]=8'b11111111;
memory[11248]=8'b11111111;
memory[11249]=8'b11011111;
memory[11250]=8'b11001111;
memory[11251]=8'b00111111;
memory[11252]=8'b11000000;
memory[11253]=8'b00000000;
memory[11254]=8'b00011111;
memory[11255]=8'b11111000;
memory[11256]=8'b00000000;
memory[11257]=8'b00000000;
memory[11258]=8'b00111111;
memory[11259]=8'b11111111;
memory[11260]=8'b00000000;
memory[11261]=8'b01111111;
memory[11262]=8'b11111111;
memory[11263]=8'b11111111;
memory[11264]=8'b10000000;
memory[11265]=8'b00111111;
memory[11266]=8'b11111111;
memory[11267]=8'b11111111;
memory[11268]=8'b11011111;
memory[11269]=8'b11111111;
memory[11270]=8'b11111111;
memory[11271]=8'b11111111;
memory[11272]=8'b11111111;
memory[11273]=8'b11111111;
memory[11274]=8'b11111111;
memory[11275]=8'b11111111;
memory[11276]=8'b11111111;
memory[11277]=8'b11111111;
memory[11278]=8'b11111111;
memory[11279]=8'b11111111;
memory[11280]=8'b11111111;
memory[11281]=8'b11111111;
memory[11282]=8'b11111111;
memory[11283]=8'b11111111;
memory[11284]=8'b11111111;
memory[11285]=8'b11111111;
memory[11286]=8'b11111111;
memory[11287]=8'b11111111;
memory[11288]=8'b11111111;
memory[11289]=8'b00011111;
memory[11290]=8'b10011110;
memory[11291]=8'b00111110;
memory[11292]=8'b00000000;
memory[11293]=8'b00000000;
memory[11294]=8'b00000111;
memory[11295]=8'b11100000;
memory[11296]=8'b00000000;
memory[11297]=8'b00000000;
memory[11298]=8'b00011111;
memory[11299]=8'b11111110;
memory[11300]=8'b00000000;
memory[11301]=8'b01111100;
memory[11302]=8'b11111111;
memory[11303]=8'b11111111;
memory[11304]=8'b11000000;
memory[11305]=8'b00111111;
memory[11306]=8'b11111111;
memory[11307]=8'b11111111;
memory[11308]=8'b11111111;
memory[11309]=8'b11111111;
memory[11310]=8'b11111111;
memory[11311]=8'b11111111;
memory[11312]=8'b11111111;
memory[11313]=8'b11111111;
memory[11314]=8'b11111111;
memory[11315]=8'b11111111;
memory[11316]=8'b11111111;
memory[11317]=8'b11111111;
memory[11318]=8'b11111111;
memory[11319]=8'b11111111;
memory[11320]=8'b11111111;
memory[11321]=8'b11111111;
memory[11322]=8'b11111111;
memory[11323]=8'b11111111;
memory[11324]=8'b11111111;
memory[11325]=8'b11111111;
memory[11326]=8'b11111111;
memory[11327]=8'b11111111;
memory[11328]=8'b11111110;
memory[11329]=8'b00111111;
memory[11330]=8'b10001100;
memory[11331]=8'b01111100;
memory[11332]=8'b00000000;
memory[11333]=8'b00000000;
memory[11334]=8'b00001111;
memory[11335]=8'b11100000;
memory[11336]=8'b00000000;
memory[11337]=8'b00000000;
memory[11338]=8'b00011111;
memory[11339]=8'b11111110;
memory[11340]=8'b00000000;
memory[11341]=8'b01111000;
memory[11342]=8'b00111111;
memory[11343]=8'b11111111;
memory[11344]=8'b11000000;
memory[11345]=8'b00111111;
memory[11346]=8'b11111111;
memory[11347]=8'b11111111;
memory[11348]=8'b11111111;
memory[11349]=8'b11111111;
memory[11350]=8'b11111111;
memory[11351]=8'b11111111;
memory[11352]=8'b11111111;
memory[11353]=8'b11111111;
memory[11354]=8'b11111111;
memory[11355]=8'b11111111;
memory[11356]=8'b11111111;
memory[11357]=8'b11111111;
memory[11358]=8'b11111111;
memory[11359]=8'b11111111;
memory[11360]=8'b11111111;
memory[11361]=8'b11111111;
memory[11362]=8'b11111111;
memory[11363]=8'b11111111;
memory[11364]=8'b11111111;
memory[11365]=8'b11111111;
memory[11366]=8'b11111111;
memory[11367]=8'b11111111;
memory[11368]=8'b11111100;
memory[11369]=8'b00011111;
memory[11370]=8'b10000000;
memory[11371]=8'b01111000;
memory[11372]=8'b00000000;
memory[11373]=8'b00000000;
memory[11374]=8'b00011111;
memory[11375]=8'b11100000;
memory[11376]=8'b00000000;
memory[11377]=8'b00000000;
memory[11378]=8'b00001111;
memory[11379]=8'b11111110;
memory[11380]=8'b00000000;
memory[11381]=8'b01111000;
memory[11382]=8'b00111111;
memory[11383]=8'b11111111;
memory[11384]=8'b11000000;
memory[11385]=8'b00111111;
memory[11386]=8'b11111111;
memory[11387]=8'b11111111;
memory[11388]=8'b11111111;
memory[11389]=8'b11111111;
memory[11390]=8'b11111111;
memory[11391]=8'b11111111;
memory[11392]=8'b11111111;
memory[11393]=8'b11111111;
memory[11394]=8'b11111111;
memory[11395]=8'b11111111;
memory[11396]=8'b11111111;
memory[11397]=8'b11111111;
memory[11398]=8'b11111111;
memory[11399]=8'b11111111;
memory[11400]=8'b11111111;
memory[11401]=8'b11111111;
memory[11402]=8'b11111111;
memory[11403]=8'b11111111;
memory[11404]=8'b11111111;
memory[11405]=8'b11111111;
memory[11406]=8'b11111111;
memory[11407]=8'b11111111;
memory[11408]=8'b11110000;
memory[11409]=8'b00000111;
memory[11410]=8'b10000000;
memory[11411]=8'b00110000;
memory[11412]=8'b00000000;
memory[11413]=8'b00000001;
memory[11414]=8'b11111111;
memory[11415]=8'b11100000;
memory[11416]=8'b00000000;
memory[11417]=8'b00000000;
memory[11418]=8'b00001111;
memory[11419]=8'b11111100;
memory[11420]=8'b00000000;
memory[11421]=8'b01111100;
memory[11422]=8'b01111111;
memory[11423]=8'b11111111;
memory[11424]=8'b11000000;
memory[11425]=8'b01111111;
memory[11426]=8'b11111111;
memory[11427]=8'b11111111;
memory[11428]=8'b11111111;
memory[11429]=8'b11111111;
memory[11430]=8'b11111111;
memory[11431]=8'b11111111;
memory[11432]=8'b11111111;
memory[11433]=8'b11111111;
memory[11434]=8'b11111111;
memory[11435]=8'b11111111;
memory[11436]=8'b11111111;
memory[11437]=8'b11111111;
memory[11438]=8'b11111111;
memory[11439]=8'b11111111;
memory[11440]=8'b11111111;
memory[11441]=8'b11111111;
memory[11442]=8'b11111111;
memory[11443]=8'b11111111;
memory[11444]=8'b11111111;
memory[11445]=8'b11111111;
memory[11446]=8'b11111111;
memory[11447]=8'b11111111;
memory[11448]=8'b11100000;
memory[11449]=8'b00000110;
memory[11450]=8'b00000000;
memory[11451]=8'b00000000;
memory[11452]=8'b00000000;
memory[11453]=8'b00001111;
memory[11454]=8'b11111111;
memory[11455]=8'b11100000;
memory[11456]=8'b00000000;
memory[11457]=8'b00000000;
memory[11458]=8'b00001111;
memory[11459]=8'b11111100;
memory[11460]=8'b00000000;
memory[11461]=8'b00111100;
memory[11462]=8'b01111111;
memory[11463]=8'b11111111;
memory[11464]=8'b10000000;
memory[11465]=8'b01111111;
memory[11466]=8'b11111111;
memory[11467]=8'b11111111;
memory[11468]=8'b11111111;
memory[11469]=8'b11111111;
memory[11470]=8'b11111111;
memory[11471]=8'b11111111;
memory[11472]=8'b11111111;
memory[11473]=8'b11111111;
memory[11474]=8'b11111111;
memory[11475]=8'b11111111;
memory[11476]=8'b11111111;
memory[11477]=8'b11111111;
memory[11478]=8'b11111111;
memory[11479]=8'b11111111;
memory[11480]=8'b11111111;
memory[11481]=8'b11111111;
memory[11482]=8'b11111111;
memory[11483]=8'b11111111;
memory[11484]=8'b11111111;
memory[11485]=8'b11111111;
memory[11486]=8'b11111111;
memory[11487]=8'b11111111;
memory[11488]=8'b10000000;
memory[11489]=8'b00000000;
memory[11490]=8'b00000000;
memory[11491]=8'b00000000;
memory[11492]=8'b00000001;
memory[11493]=8'b11111111;
memory[11494]=8'b11100000;
memory[11495]=8'b00000000;
memory[11496]=8'b00000000;
memory[11497]=8'b00000000;
memory[11498]=8'b00000011;
memory[11499]=8'b11110000;
memory[11500]=8'b00000000;
memory[11501]=8'b00111100;
memory[11502]=8'b11111111;
memory[11503]=8'b11111111;
memory[11504]=8'b00000000;
memory[11505]=8'b01111111;
memory[11506]=8'b11111111;
memory[11507]=8'b11111111;
memory[11508]=8'b11111111;
memory[11509]=8'b11111111;
memory[11510]=8'b11111111;
memory[11511]=8'b11111111;
memory[11512]=8'b11111111;
memory[11513]=8'b11111111;
memory[11514]=8'b11111111;
memory[11515]=8'b11111111;
memory[11516]=8'b11111111;
memory[11517]=8'b11111111;
memory[11518]=8'b11111111;
memory[11519]=8'b11111111;
memory[11520]=8'b11111111;
memory[11521]=8'b11111111;
memory[11522]=8'b11111111;
memory[11523]=8'b11111111;
memory[11524]=8'b11111111;
memory[11525]=8'b11111111;
memory[11526]=8'b11111111;
memory[11527]=8'b11111110;
memory[11528]=8'b00000000;
memory[11529]=8'b00000000;
memory[11530]=8'b00000000;
memory[11531]=8'b00000000;
memory[11532]=8'b01111111;
memory[11533]=8'b11111111;
memory[11534]=8'b11100000;
memory[11535]=8'b00000000;
memory[11536]=8'b00000000;
memory[11537]=8'b00000000;
memory[11538]=8'b00000000;
memory[11539]=8'b00000000;
memory[11540]=8'b00000000;
memory[11541]=8'b01111111;
memory[11542]=8'b11111111;
memory[11543]=8'b11111110;
memory[11544]=8'b00000000;
memory[11545]=8'b11111111;
memory[11546]=8'b11111111;
memory[11547]=8'b11111111;
memory[11548]=8'b11111111;
memory[11549]=8'b11111111;
memory[11550]=8'b11111111;
memory[11551]=8'b11111111;
memory[11552]=8'b11111111;
memory[11553]=8'b11111111;
memory[11554]=8'b11111111;
memory[11555]=8'b11111111;
memory[11556]=8'b11111111;
memory[11557]=8'b11111111;
memory[11558]=8'b11111111;
memory[11559]=8'b11111111;
memory[11560]=8'b11111111;
memory[11561]=8'b11111111;
memory[11562]=8'b11111111;
memory[11563]=8'b11111111;
memory[11564]=8'b11111111;
memory[11565]=8'b11111111;
memory[11566]=8'b11111111;
memory[11567]=8'b11111000;
memory[11568]=8'b00000000;
memory[11569]=8'b00111000;
memory[11570]=8'b00111111;
memory[11571]=8'b11111111;
memory[11572]=8'b11111111;
memory[11573]=8'b11111111;
memory[11574]=8'b11110000;
memory[11575]=8'b00000000;
memory[11576]=8'b00000000;
memory[11577]=8'b00000000;
memory[11578]=8'b00000000;
memory[11579]=8'b00000000;
memory[11580]=8'b00000000;
memory[11581]=8'b01111111;
memory[11582]=8'b11111111;
memory[11583]=8'b11111100;
memory[11584]=8'b00000001;
memory[11585]=8'b11111111;
memory[11586]=8'b11111111;
memory[11587]=8'b11111111;
memory[11588]=8'b11111111;
memory[11589]=8'b11111111;
memory[11590]=8'b11111111;
memory[11591]=8'b11111111;
memory[11592]=8'b11111111;
memory[11593]=8'b11111111;
memory[11594]=8'b11111111;
memory[11595]=8'b11111111;
memory[11596]=8'b11111111;
memory[11597]=8'b11111111;
memory[11598]=8'b11111111;
memory[11599]=8'b11111111;
memory[11600]=8'b11111111;
memory[11601]=8'b11111111;
memory[11602]=8'b11111111;
memory[11603]=8'b11111111;
memory[11604]=8'b11111111;
memory[11605]=8'b11111111;
memory[11606]=8'b11111111;
memory[11607]=8'b11110000;
memory[11608]=8'b00000000;
memory[11609]=8'b11111001;
memory[11610]=8'b11111111;
memory[11611]=8'b11111111;
memory[11612]=8'b11111111;
memory[11613]=8'b11001111;
memory[11614]=8'b11111110;
memory[11615]=8'b00000000;
memory[11616]=8'b00000000;
memory[11617]=8'b00000000;
memory[11618]=8'b00000000;
memory[11619]=8'b00000000;
memory[11620]=8'b00000000;
memory[11621]=8'b01111111;
memory[11622]=8'b11111111;
memory[11623]=8'b11111100;
memory[11624]=8'b00000011;
memory[11625]=8'b11111111;
memory[11626]=8'b11111111;
memory[11627]=8'b11111111;
memory[11628]=8'b11111111;
memory[11629]=8'b11111111;
memory[11630]=8'b11111111;
memory[11631]=8'b11111111;
memory[11632]=8'b11111111;
memory[11633]=8'b11111111;
memory[11634]=8'b11111111;
memory[11635]=8'b11111111;
memory[11636]=8'b11111111;
memory[11637]=8'b11111111;
memory[11638]=8'b11111111;
memory[11639]=8'b11111111;
memory[11640]=8'b11111111;
memory[11641]=8'b11111111;
memory[11642]=8'b11111111;
memory[11643]=8'b11111111;
memory[11644]=8'b11111111;
memory[11645]=8'b11111111;
memory[11646]=8'b11111111;
memory[11647]=8'b11000000;
memory[11648]=8'b00000001;
memory[11649]=8'b11111111;
memory[11650]=8'b11111111;
memory[11651]=8'b11111111;
memory[11652]=8'b11111111;
memory[11653]=8'b11000011;
memory[11654]=8'b11111111;
memory[11655]=8'b00000000;
memory[11656]=8'b00000000;
memory[11657]=8'b00000000;
memory[11658]=8'b00000000;
memory[11659]=8'b00000000;
memory[11660]=8'b00000000;
memory[11661]=8'b01111111;
memory[11662]=8'b11111111;
memory[11663]=8'b11111000;
memory[11664]=8'b00000111;
memory[11665]=8'b11111111;
memory[11666]=8'b11111111;
memory[11667]=8'b11111111;
memory[11668]=8'b11111111;
memory[11669]=8'b11111111;
memory[11670]=8'b11111111;
memory[11671]=8'b11111111;
memory[11672]=8'b11111111;
memory[11673]=8'b11111111;
memory[11674]=8'b11111111;
memory[11675]=8'b11111111;
memory[11676]=8'b11111111;
memory[11677]=8'b11111111;
memory[11678]=8'b11111111;
memory[11679]=8'b11111111;
memory[11680]=8'b11111111;
memory[11681]=8'b11111111;
memory[11682]=8'b11111111;
memory[11683]=8'b11111111;
memory[11684]=8'b11111111;
memory[11685]=8'b11111111;
memory[11686]=8'b11111111;
memory[11687]=8'b11000000;
memory[11688]=8'b00000011;
memory[11689]=8'b11111111;
memory[11690]=8'b11111111;
memory[11691]=8'b11111100;
memory[11692]=8'b01111111;
memory[11693]=8'b11000000;
memory[11694]=8'b00000000;
memory[11695]=8'b00000000;
memory[11696]=8'b00000000;
memory[11697]=8'b00000000;
memory[11698]=8'b00000000;
memory[11699]=8'b00000000;
memory[11700]=8'b00000000;
memory[11701]=8'b11111111;
memory[11702]=8'b11111111;
memory[11703]=8'b11110000;
memory[11704]=8'b00001111;
memory[11705]=8'b11111111;
memory[11706]=8'b11111111;
memory[11707]=8'b11111111;
memory[11708]=8'b11111111;
memory[11709]=8'b11111111;
memory[11710]=8'b11111111;
memory[11711]=8'b11111111;
memory[11712]=8'b11111111;
memory[11713]=8'b11111111;
memory[11714]=8'b11111111;
memory[11715]=8'b11111111;
memory[11716]=8'b11111111;
memory[11717]=8'b11111111;
memory[11718]=8'b11111111;
memory[11719]=8'b11111111;
memory[11720]=8'b11111111;
memory[11721]=8'b11111111;
memory[11722]=8'b11111111;
memory[11723]=8'b11111111;
memory[11724]=8'b11111111;
memory[11725]=8'b11111111;
memory[11726]=8'b11111111;
memory[11727]=8'b11100000;
memory[11728]=8'b00000111;
memory[11729]=8'b11111111;
memory[11730]=8'b11111111;
memory[11731]=8'b11111000;
memory[11732]=8'b00000111;
memory[11733]=8'b10000000;
memory[11734]=8'b00000000;
memory[11735]=8'b00000000;
memory[11736]=8'b00000000;
memory[11737]=8'b00000000;
memory[11738]=8'b00000000;
memory[11739]=8'b00000000;
memory[11740]=8'b00000001;
memory[11741]=8'b11111111;
memory[11742]=8'b11111111;
memory[11743]=8'b11100000;
memory[11744]=8'b00011111;
memory[11745]=8'b11111111;
memory[11746]=8'b11111111;
memory[11747]=8'b11111111;
memory[11748]=8'b11111111;
memory[11749]=8'b11111111;
memory[11750]=8'b11111111;
memory[11751]=8'b11111111;
memory[11752]=8'b11111111;
memory[11753]=8'b11111111;
memory[11754]=8'b11111111;
memory[11755]=8'b11111111;
memory[11756]=8'b11111111;
memory[11757]=8'b11111111;
memory[11758]=8'b11111111;
memory[11759]=8'b11111111;
memory[11760]=8'b11111111;
memory[11761]=8'b11111111;
memory[11762]=8'b11111111;
memory[11763]=8'b11111111;
memory[11764]=8'b11111111;
memory[11765]=8'b11111111;
memory[11766]=8'b11111111;
memory[11767]=8'b11000000;
memory[11768]=8'b00011111;
memory[11769]=8'b11000000;
memory[11770]=8'b00001111;
memory[11771]=8'b11110000;
memory[11772]=8'b00000000;
memory[11773]=8'b00000000;
memory[11774]=8'b00000000;
memory[11775]=8'b00000000;
memory[11776]=8'b00000000;
memory[11777]=8'b00000000;
memory[11778]=8'b00000000;
memory[11779]=8'b00000000;
memory[11780]=8'b00000011;
memory[11781]=8'b11111111;
memory[11782]=8'b11111111;
memory[11783]=8'b11000000;
memory[11784]=8'b00111111;
memory[11785]=8'b11111111;
memory[11786]=8'b11111111;
memory[11787]=8'b11111111;
memory[11788]=8'b11111111;
memory[11789]=8'b11111111;
memory[11790]=8'b11111111;
memory[11791]=8'b11111111;
memory[11792]=8'b11111111;
memory[11793]=8'b11111111;
memory[11794]=8'b11111111;
memory[11795]=8'b11111111;
memory[11796]=8'b11111111;
memory[11797]=8'b11111111;
memory[11798]=8'b11111111;
memory[11799]=8'b11111111;
memory[11800]=8'b11111111;
memory[11801]=8'b11111111;
memory[11802]=8'b11111111;
memory[11803]=8'b11111111;
memory[11804]=8'b11111111;
memory[11805]=8'b11111111;
memory[11806]=8'b11111111;
memory[11807]=8'b10000001;
memory[11808]=8'b11111110;
memory[11809]=8'b00000000;
memory[11810]=8'b00000000;
memory[11811]=8'b00000000;
memory[11812]=8'b00000000;
memory[11813]=8'b00000000;
memory[11814]=8'b00000000;
memory[11815]=8'b00000001;
memory[11816]=8'b11111000;
memory[11817]=8'b00000000;
memory[11818]=8'b00000000;
memory[11819]=8'b00000000;
memory[11820]=8'b00000111;
memory[11821]=8'b11111111;
memory[11822]=8'b11111111;
memory[11823]=8'b00000000;
memory[11824]=8'b11111111;
memory[11825]=8'b11111111;
memory[11826]=8'b11111111;
memory[11827]=8'b11111111;
memory[11828]=8'b11111111;
memory[11829]=8'b11111111;
memory[11830]=8'b11111111;
memory[11831]=8'b11111111;
memory[11832]=8'b11111111;
memory[11833]=8'b11111111;
memory[11834]=8'b11111111;
memory[11835]=8'b11111111;
memory[11836]=8'b11111111;
memory[11837]=8'b11111111;
memory[11838]=8'b11111111;
memory[11839]=8'b11111111;
memory[11840]=8'b11111111;
memory[11841]=8'b11111111;
memory[11842]=8'b11111111;
memory[11843]=8'b11111111;
memory[11844]=8'b11111111;
memory[11845]=8'b11111111;
memory[11846]=8'b11111111;
memory[11847]=8'b00001111;
memory[11848]=8'b11110000;
memory[11849]=8'b00000111;
memory[11850]=8'b11111000;
memory[11851]=8'b00000000;
memory[11852]=8'b00000000;
memory[11853]=8'b00000000;
memory[11854]=8'b00000000;
memory[11855]=8'b00111111;
memory[11856]=8'b11111111;
memory[11857]=8'b10000000;
memory[11858]=8'b00000000;
memory[11859]=8'b00000000;
memory[11860]=8'b00111111;
memory[11861]=8'b11111111;
memory[11862]=8'b11111110;
memory[11863]=8'b00000001;
memory[11864]=8'b11111111;
memory[11865]=8'b11111111;
memory[11866]=8'b11111111;
memory[11867]=8'b11111111;
memory[11868]=8'b11111111;
memory[11869]=8'b11111111;
memory[11870]=8'b11111111;
memory[11871]=8'b11111111;
memory[11872]=8'b11111111;
memory[11873]=8'b11111111;
memory[11874]=8'b11111111;
memory[11875]=8'b11111111;
memory[11876]=8'b11111111;
memory[11877]=8'b11111111;
memory[11878]=8'b11111111;
memory[11879]=8'b11111111;
memory[11880]=8'b11111111;
memory[11881]=8'b11111111;
memory[11882]=8'b11111111;
memory[11883]=8'b11111111;
memory[11884]=8'b11111111;
memory[11885]=8'b11111111;
memory[11886]=8'b11111111;
memory[11887]=8'b11111111;
memory[11888]=8'b10000000;
memory[11889]=8'b00111111;
memory[11890]=8'b11111111;
memory[11891]=8'b11100000;
memory[11892]=8'b00000000;
memory[11893]=8'b00000000;
memory[11894]=8'b00000001;
memory[11895]=8'b11111111;
memory[11896]=8'b11111111;
memory[11897]=8'b11111100;
memory[11898]=8'b00000000;
memory[11899]=8'b00000001;
memory[11900]=8'b11111111;
memory[11901]=8'b11111111;
memory[11902]=8'b11111110;
memory[11903]=8'b00000011;
memory[11904]=8'b11111111;
memory[11905]=8'b11111111;
memory[11906]=8'b11111111;
memory[11907]=8'b11111111;
memory[11908]=8'b11111111;
memory[11909]=8'b11111111;
memory[11910]=8'b11111111;
memory[11911]=8'b11111111;
memory[11912]=8'b11111111;
memory[11913]=8'b11111111;
memory[11914]=8'b11111111;
memory[11915]=8'b11111111;
memory[11916]=8'b11111111;
memory[11917]=8'b11111111;
memory[11918]=8'b11111111;
memory[11919]=8'b11111111;
memory[11920]=8'b11111111;
memory[11921]=8'b11111111;
memory[11922]=8'b11111111;
memory[11923]=8'b11111111;
memory[11924]=8'b11111111;
memory[11925]=8'b11111111;
memory[11926]=8'b11111111;
memory[11927]=8'b11111110;
memory[11928]=8'b00000000;
memory[11929]=8'b11111100;
memory[11930]=8'b11111111;
memory[11931]=8'b11111111;
memory[11932]=8'b00000000;
memory[11933]=8'b00000000;
memory[11934]=8'b00011111;
memory[11935]=8'b11111000;
memory[11936]=8'b00000001;
memory[11937]=8'b11111111;
memory[11938]=8'b11100000;
memory[11939]=8'b00111111;
memory[11940]=8'b11111111;
memory[11941]=8'b11111111;
memory[11942]=8'b11111100;
memory[11943]=8'b00000111;
memory[11944]=8'b11111111;
memory[11945]=8'b11111111;
memory[11946]=8'b11111111;
memory[11947]=8'b11111111;
memory[11948]=8'b11111111;
memory[11949]=8'b11111111;
memory[11950]=8'b11111111;
memory[11951]=8'b11111111;
memory[11952]=8'b11111111;
memory[11953]=8'b11111111;
memory[11954]=8'b11111111;
memory[11955]=8'b11111111;
memory[11956]=8'b11111111;
memory[11957]=8'b11111111;
memory[11958]=8'b11111111;
memory[11959]=8'b11111111;
memory[11960]=8'b11111111;
memory[11961]=8'b11111111;
memory[11962]=8'b11111111;
memory[11963]=8'b11111111;
memory[11964]=8'b11111111;
memory[11965]=8'b11111111;
memory[11966]=8'b11111111;
memory[11967]=8'b11111000;
memory[11968]=8'b00000001;
memory[11969]=8'b11111110;
memory[11970]=8'b00000000;
memory[11971]=8'b11111111;
memory[11972]=8'b11111100;
memory[11973]=8'b00000001;
memory[11974]=8'b11111111;
memory[11975]=8'b00000000;
memory[11976]=8'b01110000;
memory[11977]=8'b00001111;
memory[11978]=8'b11111111;
memory[11979]=8'b11111111;
memory[11980]=8'b11111111;
memory[11981]=8'b11111111;
memory[11982]=8'b11111000;
memory[11983]=8'b00001111;
memory[11984]=8'b11111111;
memory[11985]=8'b11111111;
memory[11986]=8'b00000000;
memory[11987]=8'b00000000;
memory[11988]=8'b01111111;
memory[11989]=8'b11111111;
memory[11990]=8'b11111111;
memory[11991]=8'b11111111;
memory[11992]=8'b11111111;
memory[11993]=8'b11111111;
memory[11994]=8'b11111111;
memory[11995]=8'b11111111;
memory[11996]=8'b11111111;
memory[11997]=8'b11111111;
memory[11998]=8'b11111111;
memory[11999]=8'b11111111;
memory[12000]=8'b11111111;
memory[12001]=8'b11111111;
memory[12002]=8'b11111111;
memory[12003]=8'b11111111;
memory[12004]=8'b11111111;
memory[12005]=8'b11111111;
memory[12006]=8'b11111111;
memory[12007]=8'b11110000;
memory[12008]=8'b00000011;
memory[12009]=8'b11111111;
memory[12010]=8'b11111111;
memory[12011]=8'b10000111;
memory[12012]=8'b11111111;
memory[12013]=8'b11111111;
memory[12014]=8'b11111000;
memory[12015]=8'b00011111;
memory[12016]=8'b11111111;
memory[12017]=8'b11111111;
memory[12018]=8'b11111111;
memory[12019]=8'b11111111;
memory[12020]=8'b11111111;
memory[12021]=8'b11111111;
memory[12022]=8'b11110000;
memory[12023]=8'b00011111;
memory[12024]=8'b11111111;
memory[12025]=8'b11110000;
memory[12026]=8'b00000001;
memory[12027]=8'b11111111;
memory[12028]=8'b11111111;
memory[12029]=8'b11111111;
memory[12030]=8'b11111111;
memory[12031]=8'b11111111;
memory[12032]=8'b11111111;
memory[12033]=8'b11111111;
memory[12034]=8'b11111111;
memory[12035]=8'b11111111;
memory[12036]=8'b11111111;
memory[12037]=8'b11111111;
memory[12038]=8'b11111111;
memory[12039]=8'b11111111;
memory[12040]=8'b11111111;
memory[12041]=8'b11111111;
memory[12042]=8'b11111111;
memory[12043]=8'b11111111;
memory[12044]=8'b11111111;
memory[12045]=8'b11111111;
memory[12046]=8'b11111111;
memory[12047]=8'b11100000;
memory[12048]=8'b00001111;
memory[12049]=8'b11111111;
memory[12050]=8'b11111111;
memory[12051]=8'b11111000;
memory[12052]=8'b00000011;
memory[12053]=8'b11111111;
memory[12054]=8'b00000000;
memory[12055]=8'b11111111;
memory[12056]=8'b11111111;
memory[12057]=8'b11111111;
memory[12058]=8'b11111111;
memory[12059]=8'b11111111;
memory[12060]=8'b11111111;
memory[12061]=8'b11111111;
memory[12062]=8'b11100000;
memory[12063]=8'b00111111;
memory[12064]=8'b11111111;
memory[12065]=8'b11000000;
memory[12066]=8'b00000011;
memory[12067]=8'b11111111;
memory[12068]=8'b11111110;
memory[12069]=8'b00111111;
memory[12070]=8'b11111111;
memory[12071]=8'b11111111;
memory[12072]=8'b11111111;
memory[12073]=8'b11111111;
memory[12074]=8'b11111111;
memory[12075]=8'b11111111;
memory[12076]=8'b11111111;
memory[12077]=8'b11111111;
memory[12078]=8'b11111111;
memory[12079]=8'b11111111;
memory[12080]=8'b11111111;
memory[12081]=8'b11111111;
memory[12082]=8'b11111111;
memory[12083]=8'b11111111;
memory[12084]=8'b11111111;
memory[12085]=8'b11111111;
memory[12086]=8'b11111111;
memory[12087]=8'b11000000;
memory[12088]=8'b00111111;
memory[12089]=8'b11111111;
memory[12090]=8'b11111111;
memory[12091]=8'b11111111;
memory[12092]=8'b10000000;
memory[12093]=8'b00000000;
memory[12094]=8'b00000011;
memory[12095]=8'b11111111;
memory[12096]=8'b11111111;
memory[12097]=8'b11111111;
memory[12098]=8'b11111111;
memory[12099]=8'b11111111;
memory[12100]=8'b11111111;
memory[12101]=8'b11111111;
memory[12102]=8'b11100000;
memory[12103]=8'b00111111;
memory[12104]=8'b11111111;
memory[12105]=8'b00000000;
memory[12106]=8'b00001111;
memory[12107]=8'b11111111;
memory[12108]=8'b11111111;
memory[12109]=8'b11000111;
memory[12110]=8'b11111111;
memory[12111]=8'b11111111;
memory[12112]=8'b11111111;
memory[12113]=8'b11111111;
memory[12114]=8'b11111111;
memory[12115]=8'b11111111;
memory[12116]=8'b11111111;
memory[12117]=8'b11111111;
memory[12118]=8'b11111111;
memory[12119]=8'b11111111;
memory[12120]=8'b11111111;
memory[12121]=8'b11111111;
memory[12122]=8'b11111111;
memory[12123]=8'b11111111;
memory[12124]=8'b11111111;
memory[12125]=8'b11111111;
memory[12126]=8'b11111111;
memory[12127]=8'b10000000;
memory[12128]=8'b11111111;
memory[12129]=8'b11111111;
memory[12130]=8'b11111111;
memory[12131]=8'b11111111;
memory[12132]=8'b11110000;
memory[12133]=8'b11111100;
memory[12134]=8'b00000111;
memory[12135]=8'b11111111;
memory[12136]=8'b11111111;
memory[12137]=8'b11111111;
memory[12138]=8'b11111111;
memory[12139]=8'b11111111;
memory[12140]=8'b11111111;
memory[12141]=8'b11111111;
memory[12142]=8'b11000000;
memory[12143]=8'b01111111;
memory[12144]=8'b11111100;
memory[12145]=8'b00000000;
memory[12146]=8'b00111111;
memory[12147]=8'b11111111;
memory[12148]=8'b11111111;
memory[12149]=8'b11110000;
memory[12150]=8'b11111111;
memory[12151]=8'b11111111;
memory[12152]=8'b11111111;
memory[12153]=8'b11111111;
memory[12154]=8'b11111111;
memory[12155]=8'b11111111;
memory[12156]=8'b11111111;
memory[12157]=8'b11111111;
memory[12158]=8'b11111111;
memory[12159]=8'b11111111;
memory[12160]=8'b11111111;
memory[12161]=8'b11111111;
memory[12162]=8'b11111111;
memory[12163]=8'b11111111;
memory[12164]=8'b11111111;
memory[12165]=8'b11111111;
memory[12166]=8'b11111111;
memory[12167]=8'b11111011;
memory[12168]=8'b11111111;
memory[12169]=8'b11111111;
memory[12170]=8'b11111111;
memory[12171]=8'b11111111;
memory[12172]=8'b11110000;
memory[12173]=8'b00111110;
memory[12174]=8'b00000111;
memory[12175]=8'b11111111;
memory[12176]=8'b11111111;
memory[12177]=8'b11111111;
memory[12178]=8'b11111111;
memory[12179]=8'b11111111;
memory[12180]=8'b11111111;
memory[12181]=8'b11111111;
memory[12182]=8'b10000000;
memory[12183]=8'b11111111;
memory[12184]=8'b11111000;
memory[12185]=8'b00000000;
memory[12186]=8'b01111111;
memory[12187]=8'b11111110;
memory[12188]=8'b01111111;
memory[12189]=8'b11111110;
memory[12190]=8'b00111111;
memory[12191]=8'b11111111;
memory[12192]=8'b11111111;
memory[12193]=8'b11111111;
memory[12194]=8'b11111111;
memory[12195]=8'b11111111;
memory[12196]=8'b11111111;
memory[12197]=8'b11111111;
memory[12198]=8'b11111111;
memory[12199]=8'b11111111;
memory[12200]=8'b11111111;
memory[12201]=8'b11111111;
memory[12202]=8'b11111111;
memory[12203]=8'b11111111;
memory[12204]=8'b11111111;
memory[12205]=8'b11111111;
memory[12206]=8'b11111111;
memory[12207]=8'b11111111;
memory[12208]=8'b11111111;
memory[12209]=8'b11111111;
memory[12210]=8'b11111111;
memory[12211]=8'b11111111;
memory[12212]=8'b11111000;
memory[12213]=8'b00111110;
memory[12214]=8'b00001111;
memory[12215]=8'b11111111;
memory[12216]=8'b11111111;
memory[12217]=8'b11111111;
memory[12218]=8'b11111111;
memory[12219]=8'b11111111;
memory[12220]=8'b11111111;
memory[12221]=8'b11111111;
memory[12222]=8'b10000000;
memory[12223]=8'b11111111;
memory[12224]=8'b11110000;
memory[12225]=8'b00000000;
memory[12226]=8'b01111111;
memory[12227]=8'b11001110;
memory[12228]=8'b01111111;
memory[12229]=8'b11111111;
memory[12230]=8'b11001111;
memory[12231]=8'b11111111;
memory[12232]=8'b11111111;
memory[12233]=8'b11111111;
memory[12234]=8'b11111111;
memory[12235]=8'b11111111;
memory[12236]=8'b11111111;
memory[12237]=8'b11111111;
memory[12238]=8'b11111111;
memory[12239]=8'b11111111;
memory[12240]=8'b11111111;
memory[12241]=8'b11111111;
memory[12242]=8'b11111111;
memory[12243]=8'b11111111;
memory[12244]=8'b11111111;
memory[12245]=8'b11111111;
memory[12246]=8'b11111111;
memory[12247]=8'b11111111;
memory[12248]=8'b11111111;
memory[12249]=8'b11111111;
memory[12250]=8'b11111111;
memory[12251]=8'b11111111;
memory[12252]=8'b11111000;
memory[12253]=8'b01111110;
memory[12254]=8'b00011111;
memory[12255]=8'b11111111;
memory[12256]=8'b11111111;
memory[12257]=8'b11111111;
memory[12258]=8'b11111111;
memory[12259]=8'b11111111;
memory[12260]=8'b11111111;
memory[12261]=8'b11111111;
memory[12262]=8'b10000000;
memory[12263]=8'b11111111;
memory[12264]=8'b11100000;
memory[12265]=8'b00000000;
memory[12266]=8'b00011111;
memory[12267]=8'b11100000;
memory[12268]=8'b01111111;
memory[12269]=8'b11011111;
memory[12270]=8'b11111111;
memory[12271]=8'b11111111;
memory[12272]=8'b11111111;
memory[12273]=8'b11111111;
memory[12274]=8'b11111111;
memory[12275]=8'b11111111;
memory[12276]=8'b11111111;
memory[12277]=8'b11111111;
memory[12278]=8'b11111111;
memory[12279]=8'b11111111;
memory[12280]=8'b11111111;
memory[12281]=8'b11111111;
memory[12282]=8'b11111111;
memory[12283]=8'b11111111;
memory[12284]=8'b11111111;
memory[12285]=8'b11111111;
memory[12286]=8'b11111111;
memory[12287]=8'b11111111;
memory[12288]=8'b11111111;
memory[12289]=8'b11111111;
memory[12290]=8'b11111111;
memory[12291]=8'b11111111;
memory[12292]=8'b11111000;
memory[12293]=8'b01111100;
memory[12294]=8'b00011111;
memory[12295]=8'b11111111;
memory[12296]=8'b11111111;
memory[12297]=8'b11111111;
memory[12298]=8'b11111111;
memory[12299]=8'b11111111;
memory[12300]=8'b11111111;
memory[12301]=8'b11111111;
memory[12302]=8'b00000000;
memory[12303]=8'b11111111;
memory[12304]=8'b11100000;
memory[12305]=8'b00000001;
memory[12306]=8'b11111111;
memory[12307]=8'b11000000;
memory[12308]=8'b01111111;
memory[12309]=8'b11100111;
memory[12310]=8'b11111111;
memory[12311]=8'b11111111;
memory[12312]=8'b11111111;
memory[12313]=8'b11111111;
memory[12314]=8'b11111111;
memory[12315]=8'b11111111;
memory[12316]=8'b11111111;
memory[12317]=8'b11111111;
memory[12318]=8'b11111111;
memory[12319]=8'b11111111;
memory[12320]=8'b11111111;
memory[12321]=8'b11111111;
memory[12322]=8'b11111111;
memory[12323]=8'b11111111;
memory[12324]=8'b11111111;
memory[12325]=8'b11111111;
memory[12326]=8'b11111111;
memory[12327]=8'b11111111;
memory[12328]=8'b11111111;
memory[12329]=8'b11111111;
memory[12330]=8'b11111111;
memory[12331]=8'b11111111;
memory[12332]=8'b11111000;
memory[12333]=8'b01111100;
memory[12334]=8'b00011111;
memory[12335]=8'b11111111;
memory[12336]=8'b11111111;
memory[12337]=8'b11111111;
memory[12338]=8'b11111111;
memory[12339]=8'b11111111;
memory[12340]=8'b11111111;
memory[12341]=8'b11111111;
memory[12342]=8'b00000001;
memory[12343]=8'b11111111;
memory[12344]=8'b11000000;
memory[12345]=8'b00000000;
memory[12346]=8'b11111111;
memory[12347]=8'b10000000;
memory[12348]=8'b00000111;
memory[12349]=8'b11110011;
memory[12350]=8'b10111111;
memory[12351]=8'b11111111;
memory[12352]=8'b11111111;
memory[12353]=8'b11111111;
memory[12354]=8'b11111111;
memory[12355]=8'b11111111;
memory[12356]=8'b11111111;
memory[12357]=8'b11111111;
memory[12358]=8'b11111111;
memory[12359]=8'b11111111;
memory[12360]=8'b11111111;
memory[12361]=8'b11111111;
memory[12362]=8'b11111111;
memory[12363]=8'b11111111;
memory[12364]=8'b11111111;
memory[12365]=8'b11111111;
memory[12366]=8'b11111111;
memory[12367]=8'b11111111;
memory[12368]=8'b11111111;
memory[12369]=8'b11111111;
memory[12370]=8'b11111111;
memory[12371]=8'b11111111;
memory[12372]=8'b11111000;
memory[12373]=8'b01111100;
memory[12374]=8'b00111111;
memory[12375]=8'b11111111;
memory[12376]=8'b11111111;
memory[12377]=8'b11111111;
memory[12378]=8'b11111111;
memory[12379]=8'b11111111;
memory[12380]=8'b11111111;
memory[12381]=8'b11111111;
memory[12382]=8'b00000001;
memory[12383]=8'b11111111;
memory[12384]=8'b10000000;
memory[12385]=8'b00000000;
memory[12386]=8'b00111111;
memory[12387]=8'b00000000;
memory[12388]=8'b00000000;
memory[12389]=8'b11110011;
memory[12390]=8'b10011111;
memory[12391]=8'b01111111;
memory[12392]=8'b11111111;
memory[12393]=8'b11111111;
memory[12394]=8'b11111111;
memory[12395]=8'b11111111;
memory[12396]=8'b11111111;
memory[12397]=8'b11111111;
memory[12398]=8'b11111111;
memory[12399]=8'b11111111;
memory[12400]=8'b11111111;
memory[12401]=8'b11111111;
memory[12402]=8'b11111111;
memory[12403]=8'b11111111;
memory[12404]=8'b11111111;
memory[12405]=8'b11111111;
memory[12406]=8'b11111111;
memory[12407]=8'b11111111;
memory[12408]=8'b11111111;
memory[12409]=8'b11111111;
memory[12410]=8'b11111111;
memory[12411]=8'b11111111;
memory[12412]=8'b11111000;
memory[12413]=8'b01111000;
memory[12414]=8'b00111111;
memory[12415]=8'b11111111;
memory[12416]=8'b11111111;
memory[12417]=8'b11111111;
memory[12418]=8'b11111111;
memory[12419]=8'b11111111;
memory[12420]=8'b11111111;
memory[12421]=8'b11111111;
memory[12422]=8'b00000000;
memory[12423]=8'b11111111;
memory[12424]=8'b10000000;
memory[12425]=8'b00000000;
memory[12426]=8'b00011111;
memory[12427]=8'b00000000;
memory[12428]=8'b00000000;
memory[12429]=8'b01111001;
memory[12430]=8'b10011111;
memory[12431]=8'b00111111;
memory[12432]=8'b11111111;
memory[12433]=8'b11111111;
memory[12434]=8'b11111111;
memory[12435]=8'b11111111;
memory[12436]=8'b11111111;
memory[12437]=8'b11111111;
memory[12438]=8'b11111111;
memory[12439]=8'b11111111;
memory[12440]=8'b11111111;
memory[12441]=8'b11111111;
memory[12442]=8'b11111111;
memory[12443]=8'b11111111;
memory[12444]=8'b11111111;
memory[12445]=8'b11111111;
memory[12446]=8'b11111111;
memory[12447]=8'b11111111;
memory[12448]=8'b11111111;
memory[12449]=8'b11111111;
memory[12450]=8'b11111111;
memory[12451]=8'b11111111;
memory[12452]=8'b11111000;
memory[12453]=8'b11111000;
memory[12454]=8'b00111111;
memory[12455]=8'b11111111;
memory[12456]=8'b11111111;
memory[12457]=8'b11111111;
memory[12458]=8'b11111111;
memory[12459]=8'b11111111;
memory[12460]=8'b11111111;
memory[12461]=8'b11111111;
memory[12462]=8'b00000000;
memory[12463]=8'b11111111;
memory[12464]=8'b00000000;
memory[12465]=8'b00000000;
memory[12466]=8'b00011111;
memory[12467]=8'b11100000;
memory[12468]=8'b00000000;
memory[12469]=8'b00111000;
memory[12470]=8'b00011110;
memory[12471]=8'b00001111;
memory[12472]=8'b11111111;
memory[12473]=8'b11111111;
memory[12474]=8'b11111111;
memory[12475]=8'b11111111;
memory[12476]=8'b11111111;
memory[12477]=8'b11111111;
memory[12478]=8'b11111111;
memory[12479]=8'b11111111;
memory[12480]=8'b11111111;
memory[12481]=8'b11111111;
memory[12482]=8'b11111111;
memory[12483]=8'b11111111;
memory[12484]=8'b11111111;
memory[12485]=8'b11111111;
memory[12486]=8'b11111111;
memory[12487]=8'b11111111;
memory[12488]=8'b11111111;
memory[12489]=8'b11111111;
memory[12490]=8'b11111111;
memory[12491]=8'b11111111;
memory[12492]=8'b11111000;
memory[12493]=8'b11111000;
memory[12494]=8'b00111111;
memory[12495]=8'b11111111;
memory[12496]=8'b11111111;
memory[12497]=8'b11111111;
memory[12498]=8'b11111111;
memory[12499]=8'b11111111;
memory[12500]=8'b11111111;
memory[12501]=8'b11111111;
memory[12502]=8'b00000000;
memory[12503]=8'b01111111;
memory[12504]=8'b00000000;
memory[12505]=8'b00000000;
memory[12506]=8'b00011111;
memory[12507]=8'b11111100;
memory[12508]=8'b00000000;
memory[12509]=8'b00000000;
memory[12510]=8'b00001100;
memory[12511]=8'b00000111;
memory[12512]=8'b11111111;
memory[12513]=8'b11111111;
memory[12514]=8'b11111111;
memory[12515]=8'b11111111;
memory[12516]=8'b11111111;
memory[12517]=8'b11111111;
memory[12518]=8'b11111111;
memory[12519]=8'b11111111;
memory[12520]=8'b11111111;
memory[12521]=8'b11111111;
memory[12522]=8'b11111111;
memory[12523]=8'b11111111;
memory[12524]=8'b11111111;
memory[12525]=8'b11111111;
memory[12526]=8'b11111111;
memory[12527]=8'b11111111;
memory[12528]=8'b11111111;
memory[12529]=8'b11111111;
memory[12530]=8'b11111111;
memory[12531]=8'b11111111;
memory[12532]=8'b11111000;
memory[12533]=8'b11111000;
memory[12534]=8'b01111111;
memory[12535]=8'b11111111;
memory[12536]=8'b11111111;
memory[12537]=8'b11111111;
memory[12538]=8'b11111111;
memory[12539]=8'b11111111;
memory[12540]=8'b11111111;
memory[12541]=8'b11111111;
memory[12542]=8'b00000000;
memory[12543]=8'b00111100;
memory[12544]=8'b00000000;
memory[12545]=8'b00000000;
memory[12546]=8'b00000000;
memory[12547]=8'b01111111;
memory[12548]=8'b11110000;
memory[12549]=8'b00000000;
memory[12550]=8'b00000000;
memory[12551]=8'b00000001;
memory[12552]=8'b11111111;
memory[12553]=8'b11111111;
memory[12554]=8'b11111111;
memory[12555]=8'b11111111;
memory[12556]=8'b11111111;
memory[12557]=8'b11111111;
memory[12558]=8'b11111111;
memory[12559]=8'b11111111;
memory[12560]=8'b11111111;
memory[12561]=8'b11111111;
memory[12562]=8'b11111111;
memory[12563]=8'b11111111;
memory[12564]=8'b11111111;
memory[12565]=8'b11111111;
memory[12566]=8'b11111111;
memory[12567]=8'b11111111;
memory[12568]=8'b11111111;
memory[12569]=8'b11111111;
memory[12570]=8'b11111111;
memory[12571]=8'b11111111;
memory[12572]=8'b11111000;
memory[12573]=8'b11111000;
memory[12574]=8'b01111111;
memory[12575]=8'b11111111;
memory[12576]=8'b11111111;
memory[12577]=8'b11111111;
memory[12578]=8'b11111111;
memory[12579]=8'b11111111;
memory[12580]=8'b11111111;
memory[12581]=8'b11111111;
memory[12582]=8'b00000000;
memory[12583]=8'b00000000;
memory[12584]=8'b00000000;
memory[12585]=8'b00000000;
memory[12586]=8'b00000000;
memory[12587]=8'b01111111;
memory[12588]=8'b11111111;
memory[12589]=8'b00000000;
memory[12590]=8'b00000000;
memory[12591]=8'b00000000;
memory[12592]=8'b01111111;
memory[12593]=8'b11111111;
memory[12594]=8'b11111111;
memory[12595]=8'b11111111;
memory[12596]=8'b11111111;
memory[12597]=8'b11111111;
memory[12598]=8'b11111111;
memory[12599]=8'b11111111;
memory[12600]=8'b11111111;
memory[12601]=8'b11111111;
memory[12602]=8'b11111111;
memory[12603]=8'b11111111;
memory[12604]=8'b11111111;
memory[12605]=8'b11111111;
memory[12606]=8'b11111111;
memory[12607]=8'b11111111;
memory[12608]=8'b11111111;
memory[12609]=8'b11111111;
memory[12610]=8'b11111111;
memory[12611]=8'b11111111;
memory[12612]=8'b11111000;
memory[12613]=8'b11110000;
memory[12614]=8'b11111111;
memory[12615]=8'b11111111;
memory[12616]=8'b11111111;
memory[12617]=8'b11111111;
memory[12618]=8'b11111111;
memory[12619]=8'b11111111;
memory[12620]=8'b11111111;
memory[12621]=8'b11111111;
memory[12622]=8'b00000000;
memory[12623]=8'b00000000;
memory[12624]=8'b00000000;
memory[12625]=8'b00000000;
memory[12626]=8'b00000001;
memory[12627]=8'b11111111;
memory[12628]=8'b11111111;
memory[12629]=8'b11111111;
memory[12630]=8'b11110011;
memory[12631]=8'b11000000;
memory[12632]=8'b00011111;
memory[12633]=8'b11111111;
memory[12634]=8'b11111111;
memory[12635]=8'b11111111;
memory[12636]=8'b11111111;
memory[12637]=8'b11111111;
memory[12638]=8'b11111111;
memory[12639]=8'b11111111;
memory[12640]=8'b11111111;
memory[12641]=8'b11111111;
memory[12642]=8'b11111111;
memory[12643]=8'b11111111;
memory[12644]=8'b11111111;
memory[12645]=8'b11111111;
memory[12646]=8'b11111111;
memory[12647]=8'b11111111;
memory[12648]=8'b11111111;
memory[12649]=8'b11111111;
memory[12650]=8'b11111111;
memory[12651]=8'b11111111;
memory[12652]=8'b11110000;
memory[12653]=8'b11110000;
memory[12654]=8'b11111111;
memory[12655]=8'b11111111;
memory[12656]=8'b11111111;
memory[12657]=8'b11111111;
memory[12658]=8'b11111111;
memory[12659]=8'b11111111;
memory[12660]=8'b11111111;
memory[12661]=8'b11111111;
memory[12662]=8'b00000000;
memory[12663]=8'b00000000;
memory[12664]=8'b00000000;
memory[12665]=8'b00000000;
memory[12666]=8'b00000011;
memory[12667]=8'b11111000;
memory[12668]=8'b11111111;
memory[12669]=8'b11111111;
memory[12670]=8'b11111111;
memory[12671]=8'b11000000;
memory[12672]=8'b00001111;
memory[12673]=8'b11111111;
memory[12674]=8'b11111111;
memory[12675]=8'b11111111;
memory[12676]=8'b11111111;
memory[12677]=8'b11111111;
memory[12678]=8'b11111111;
memory[12679]=8'b11111111;
memory[12680]=8'b11111111;
memory[12681]=8'b11111111;
memory[12682]=8'b11111111;
memory[12683]=8'b11111111;
memory[12684]=8'b11111111;
memory[12685]=8'b11111111;
memory[12686]=8'b11111111;
memory[12687]=8'b11111111;
memory[12688]=8'b11111111;
memory[12689]=8'b11111111;
memory[12690]=8'b11111111;
memory[12691]=8'b11111111;
memory[12692]=8'b11110001;
memory[12693]=8'b11110000;
memory[12694]=8'b11111111;
memory[12695]=8'b11111111;
memory[12696]=8'b11111111;
memory[12697]=8'b11111111;
memory[12698]=8'b11111111;
memory[12699]=8'b11111111;
memory[12700]=8'b11111111;
memory[12701]=8'b11111111;
memory[12702]=8'b10000000;
memory[12703]=8'b00000000;
memory[12704]=8'b00000000;
memory[12705]=8'b00000000;
memory[12706]=8'b00000000;
memory[12707]=8'b00000000;
memory[12708]=8'b11111100;
memory[12709]=8'b01111111;
memory[12710]=8'b11111111;
memory[12711]=8'b11110000;
memory[12712]=8'b00001111;
memory[12713]=8'b11111111;
memory[12714]=8'b11111111;
memory[12715]=8'b11111111;
memory[12716]=8'b11111111;
memory[12717]=8'b11111111;
memory[12718]=8'b11111111;
memory[12719]=8'b11111111;
memory[12720]=8'b11111111;
memory[12721]=8'b11111111;
memory[12722]=8'b11111111;
memory[12723]=8'b11111111;
memory[12724]=8'b11111111;
memory[12725]=8'b11111111;
memory[12726]=8'b11111111;
memory[12727]=8'b11111111;
memory[12728]=8'b11111111;
memory[12729]=8'b11111111;
memory[12730]=8'b11111111;
memory[12731]=8'b11111111;
memory[12732]=8'b11110001;
memory[12733]=8'b11110001;
memory[12734]=8'b11111111;
memory[12735]=8'b11111111;
memory[12736]=8'b11111111;
memory[12737]=8'b11111111;
memory[12738]=8'b11111111;
memory[12739]=8'b11111111;
memory[12740]=8'b11111111;
memory[12741]=8'b11111111;
memory[12742]=8'b11000000;
memory[12743]=8'b00000000;
memory[12744]=8'b00000000;
memory[12745]=8'b00000000;
memory[12746]=8'b00000000;
memory[12747]=8'b00000000;
memory[12748]=8'b00000000;
memory[12749]=8'b00111111;
memory[12750]=8'b11100001;
memory[12751]=8'b11111100;
memory[12752]=8'b00001111;
memory[12753]=8'b11111111;
memory[12754]=8'b11111111;
memory[12755]=8'b11111111;
memory[12756]=8'b11111111;
memory[12757]=8'b11111111;
memory[12758]=8'b11111111;
memory[12759]=8'b11111111;
memory[12760]=8'b11111111;
memory[12761]=8'b11111111;
memory[12762]=8'b11111111;
memory[12763]=8'b11111111;
memory[12764]=8'b11111111;
memory[12765]=8'b11111111;
memory[12766]=8'b11111111;
memory[12767]=8'b11111111;
memory[12768]=8'b11111111;
memory[12769]=8'b11111111;
memory[12770]=8'b11111111;
memory[12771]=8'b11111111;
memory[12772]=8'b11110001;
memory[12773]=8'b11100001;
memory[12774]=8'b11111111;
memory[12775]=8'b11111111;
memory[12776]=8'b11111111;
memory[12777]=8'b11111111;
memory[12778]=8'b11111111;
memory[12779]=8'b11111111;
memory[12780]=8'b11111111;
memory[12781]=8'b11111111;
memory[12782]=8'b11110000;
memory[12783]=8'b00000000;
memory[12784]=8'b00000000;
memory[12785]=8'b00011111;
memory[12786]=8'b10000000;
memory[12787]=8'b00000000;
memory[12788]=8'b00000000;
memory[12789]=8'b00000000;
memory[12790]=8'b00000000;
memory[12791]=8'b00111111;
memory[12792]=8'b10000111;
memory[12793]=8'b11111111;
memory[12794]=8'b11111111;
memory[12795]=8'b11111111;
memory[12796]=8'b11111111;
memory[12797]=8'b11111111;
memory[12798]=8'b11111111;
memory[12799]=8'b11111111;
memory[12800]=8'b11111111;
memory[12801]=8'b11111111;
memory[12802]=8'b11111111;
memory[12803]=8'b11111111;
memory[12804]=8'b11111111;
memory[12805]=8'b11111111;
memory[12806]=8'b11111111;
memory[12807]=8'b11111111;
memory[12808]=8'b11111111;
memory[12809]=8'b11111111;
memory[12810]=8'b11111111;
memory[12811]=8'b11111111;
memory[12812]=8'b11110001;
memory[12813]=8'b11100001;
memory[12814]=8'b11111111;
memory[12815]=8'b11111111;
memory[12816]=8'b11111111;
memory[12817]=8'b11111111;
memory[12818]=8'b11111111;
memory[12819]=8'b11111111;
memory[12820]=8'b11111111;
memory[12821]=8'b11111111;
memory[12822]=8'b11111100;
memory[12823]=8'b00000000;
memory[12824]=8'b00000011;
memory[12825]=8'b11111111;
memory[12826]=8'b11111000;
memory[12827]=8'b00000000;
memory[12828]=8'b00000000;
memory[12829]=8'b00000111;
memory[12830]=8'b11111110;
memory[12831]=8'b00000111;
memory[12832]=8'b11110011;
memory[12833]=8'b11111111;
memory[12834]=8'b11111111;
memory[12835]=8'b11111111;
memory[12836]=8'b11111111;
memory[12837]=8'b11111111;
memory[12838]=8'b11111111;
memory[12839]=8'b11111111;
memory[12840]=8'b11111111;
memory[12841]=8'b11111111;
memory[12842]=8'b11111111;
memory[12843]=8'b11111111;
memory[12844]=8'b11111111;
memory[12845]=8'b11111111;
memory[12846]=8'b11111111;
memory[12847]=8'b11111111;
memory[12848]=8'b11111111;
memory[12849]=8'b11111111;
memory[12850]=8'b11111111;
memory[12851]=8'b11111111;
memory[12852]=8'b11100011;
memory[12853]=8'b11100001;
memory[12854]=8'b11111111;
memory[12855]=8'b11111111;
memory[12856]=8'b11111111;
memory[12857]=8'b11111111;
memory[12858]=8'b11111111;
memory[12859]=8'b11111111;
memory[12860]=8'b11111111;
memory[12861]=8'b11111111;
memory[12862]=8'b11111111;
memory[12863]=8'b11000000;
memory[12864]=8'b00111111;
memory[12865]=8'b11100000;
memory[12866]=8'b01111111;
memory[12867]=8'b10000000;
memory[12868]=8'b00000000;
memory[12869]=8'b01111111;
memory[12870]=8'b11111111;
memory[12871]=8'b10000000;
memory[12872]=8'b11111111;
memory[12873]=8'b11111111;
memory[12874]=8'b11111111;
memory[12875]=8'b11111111;
memory[12876]=8'b11111111;
memory[12877]=8'b11111111;
memory[12878]=8'b11111111;
memory[12879]=8'b11111111;
memory[12880]=8'b11111111;
memory[12881]=8'b11111111;
memory[12882]=8'b11111111;
memory[12883]=8'b11111111;
memory[12884]=8'b11111111;
memory[12885]=8'b11111111;
memory[12886]=8'b11111111;
memory[12887]=8'b11111111;
memory[12888]=8'b11111111;
memory[12889]=8'b11111111;
memory[12890]=8'b11111111;
memory[12891]=8'b11111111;
memory[12892]=8'b11100011;
memory[12893]=8'b11100001;
memory[12894]=8'b11111111;
memory[12895]=8'b11111111;
memory[12896]=8'b11111111;
memory[12897]=8'b11111111;
memory[12898]=8'b11111111;
memory[12899]=8'b11111111;
memory[12900]=8'b11111111;
memory[12901]=8'b11111111;
memory[12902]=8'b11111111;
memory[12903]=8'b11111111;
memory[12904]=8'b11111100;
memory[12905]=8'b00001100;
memory[12906]=8'b00000111;
memory[12907]=8'b11111100;
memory[12908]=8'b01111111;
memory[12909]=8'b11111000;
memory[12910]=8'b00001111;
memory[12911]=8'b11100000;
memory[12912]=8'b00111111;
memory[12913]=8'b11111111;
memory[12914]=8'b11111111;
memory[12915]=8'b11111111;
memory[12916]=8'b11111111;
memory[12917]=8'b11111111;
memory[12918]=8'b11111111;
memory[12919]=8'b11111111;
memory[12920]=8'b11111111;
memory[12921]=8'b11111111;
memory[12922]=8'b11111111;
memory[12923]=8'b11111111;
memory[12924]=8'b11111111;
memory[12925]=8'b11111111;
memory[12926]=8'b11111111;
memory[12927]=8'b11111111;
memory[12928]=8'b11111111;
memory[12929]=8'b11111111;
memory[12930]=8'b11111111;
memory[12931]=8'b11111111;
memory[12932]=8'b11100011;
memory[12933]=8'b11000001;
memory[12934]=8'b11111111;
memory[12935]=8'b11111111;
memory[12936]=8'b11111111;
memory[12937]=8'b11111111;
memory[12938]=8'b11111111;
memory[12939]=8'b11111111;
memory[12940]=8'b11111111;
memory[12941]=8'b11111111;
memory[12942]=8'b11111111;
memory[12943]=8'b11111111;
memory[12944]=8'b11111111;
memory[12945]=8'b11111111;
memory[12946]=8'b11110000;
memory[12947]=8'b11111111;
memory[12948]=8'b11111111;
memory[12949]=8'b10011111;
memory[12950]=8'b11111111;
memory[12951]=8'b11110000;
memory[12952]=8'b00011111;
memory[12953]=8'b11111111;
memory[12954]=8'b11111111;
memory[12955]=8'b11111111;
memory[12956]=8'b11111111;
memory[12957]=8'b11111111;
memory[12958]=8'b11111111;
memory[12959]=8'b11111111;
memory[12960]=8'b11111111;
memory[12961]=8'b11111111;
memory[12962]=8'b11111111;
memory[12963]=8'b11111111;
memory[12964]=8'b11111111;
memory[12965]=8'b11111111;
memory[12966]=8'b11111111;
memory[12967]=8'b11111111;
memory[12968]=8'b11111111;
memory[12969]=8'b11111111;
memory[12970]=8'b11111111;
memory[12971]=8'b11111111;
memory[12972]=8'b11100011;
memory[12973]=8'b11000001;
memory[12974]=8'b11111111;
memory[12975]=8'b11111111;
memory[12976]=8'b11111111;
memory[12977]=8'b11111111;
memory[12978]=8'b11111111;
memory[12979]=8'b11111111;
memory[12980]=8'b11111111;
memory[12981]=8'b11111111;
memory[12982]=8'b11111111;
memory[12983]=8'b11111111;
memory[12984]=8'b11111111;
memory[12985]=8'b11111111;
memory[12986]=8'b11111100;
memory[12987]=8'b00000000;
memory[12988]=8'b00000000;
memory[12989]=8'b11111111;
memory[12990]=8'b11111111;
memory[12991]=8'b11111100;
memory[12992]=8'b00001111;
memory[12993]=8'b11111111;
memory[12994]=8'b11111111;
memory[12995]=8'b11111111;
memory[12996]=8'b11111111;
memory[12997]=8'b11111111;
memory[12998]=8'b11111111;
memory[12999]=8'b11111111;
memory[13000]=8'b11111111;
memory[13001]=8'b11111111;
memory[13002]=8'b11111111;
memory[13003]=8'b11111111;
memory[13004]=8'b11111111;
memory[13005]=8'b11111111;
memory[13006]=8'b11111111;
memory[13007]=8'b11111111;
memory[13008]=8'b11111111;
memory[13009]=8'b11111111;
memory[13010]=8'b11111111;
memory[13011]=8'b11111111;
memory[13012]=8'b11100011;
memory[13013]=8'b11000011;
memory[13014]=8'b11111111;
memory[13015]=8'b11111111;
memory[13016]=8'b11111111;
memory[13017]=8'b11111111;
memory[13018]=8'b11111111;
memory[13019]=8'b11111111;
memory[13020]=8'b11111111;
memory[13021]=8'b11111111;
memory[13022]=8'b11111111;
memory[13023]=8'b11111111;
memory[13024]=8'b11111111;
memory[13025]=8'b11111111;
memory[13026]=8'b11111111;
memory[13027]=8'b00000111;
memory[13028]=8'b00001111;
memory[13029]=8'b11111111;
memory[13030]=8'b11111111;
memory[13031]=8'b11111111;
memory[13032]=8'b00000111;
memory[13033]=8'b11111111;
memory[13034]=8'b11111111;
memory[13035]=8'b11111111;
memory[13036]=8'b11111111;
memory[13037]=8'b11111111;
memory[13038]=8'b11111111;
memory[13039]=8'b11111111;
memory[13040]=8'b11111111;
memory[13041]=8'b11111111;
memory[13042]=8'b11111111;
memory[13043]=8'b11111111;
memory[13044]=8'b11111111;
memory[13045]=8'b11111111;
memory[13046]=8'b11111111;
memory[13047]=8'b11111111;
memory[13048]=8'b11111111;
memory[13049]=8'b11111111;
memory[13050]=8'b11111111;
memory[13051]=8'b11111111;
memory[13052]=8'b11100111;
memory[13053]=8'b11000011;
memory[13054]=8'b11111111;
memory[13055]=8'b11111111;
memory[13056]=8'b11111111;
memory[13057]=8'b11111111;
memory[13058]=8'b11111111;
memory[13059]=8'b11111111;
memory[13060]=8'b11111111;
memory[13061]=8'b11111111;
memory[13062]=8'b11111111;
memory[13063]=8'b11111111;
memory[13064]=8'b11111111;
memory[13065]=8'b11111111;
memory[13066]=8'b11111111;
memory[13067]=8'b00001111;
memory[13068]=8'b00001111;
memory[13069]=8'b11111111;
memory[13070]=8'b11111111;
memory[13071]=8'b11111111;
memory[13072]=8'b11111111;
memory[13073]=8'b11111111;
memory[13074]=8'b11111111;
memory[13075]=8'b11111111;
memory[13076]=8'b11111111;
memory[13077]=8'b11111111;
memory[13078]=8'b11111111;
memory[13079]=8'b11111111;
memory[13080]=8'b11111111;
memory[13081]=8'b11111111;
memory[13082]=8'b11111111;
memory[13083]=8'b11111111;
memory[13084]=8'b11111111;
memory[13085]=8'b11111111;
memory[13086]=8'b11111111;
memory[13087]=8'b11111111;
memory[13088]=8'b11111111;
memory[13089]=8'b11111111;
memory[13090]=8'b11111111;
memory[13091]=8'b11111111;
memory[13092]=8'b11000111;
memory[13093]=8'b11000011;
memory[13094]=8'b11111111;
memory[13095]=8'b11111111;
memory[13096]=8'b11111111;
memory[13097]=8'b11111111;
memory[13098]=8'b11111111;
memory[13099]=8'b11111111;
memory[13100]=8'b11111111;
memory[13101]=8'b11111111;
memory[13102]=8'b11111111;
memory[13103]=8'b11111111;
memory[13104]=8'b11111111;
memory[13105]=8'b11111111;
memory[13106]=8'b11111111;
memory[13107]=8'b10001111;
memory[13108]=8'b00001111;
memory[13109]=8'b11111111;
memory[13110]=8'b11111111;
memory[13111]=8'b11111111;
memory[13112]=8'b11111111;
memory[13113]=8'b11111111;
memory[13114]=8'b11111111;
memory[13115]=8'b11111111;
memory[13116]=8'b11111111;
memory[13117]=8'b11111111;
memory[13118]=8'b11111111;
memory[13119]=8'b11111111;
memory[13120]=8'b11111111;
memory[13121]=8'b11111111;
memory[13122]=8'b11111111;
memory[13123]=8'b11111111;
memory[13124]=8'b11111111;
memory[13125]=8'b11111111;
memory[13126]=8'b11111111;
memory[13127]=8'b11111111;
memory[13128]=8'b11111111;
memory[13129]=8'b11111111;
memory[13130]=8'b11111111;
memory[13131]=8'b11111111;
memory[13132]=8'b11000111;
memory[13133]=8'b10000111;
memory[13134]=8'b11111111;
memory[13135]=8'b11111111;
memory[13136]=8'b11111111;
memory[13137]=8'b11111111;
memory[13138]=8'b11111111;
memory[13139]=8'b11111111;
memory[13140]=8'b11111111;
memory[13141]=8'b11111111;
memory[13142]=8'b11111111;
memory[13143]=8'b11111111;
memory[13144]=8'b11111111;
memory[13145]=8'b11111111;
memory[13146]=8'b11111111;
memory[13147]=8'b10001111;
memory[13148]=8'b10001111;
memory[13149]=8'b11111111;
memory[13150]=8'b11111111;
memory[13151]=8'b11111111;
memory[13152]=8'b11111111;
memory[13153]=8'b11111111;
memory[13154]=8'b11111111;
memory[13155]=8'b11111111;
memory[13156]=8'b11111111;
memory[13157]=8'b11111111;
memory[13158]=8'b11111111;
memory[13159]=8'b11111111;
memory[13160]=8'b11111111;
memory[13161]=8'b11111111;
memory[13162]=8'b11111111;
memory[13163]=8'b11111111;
memory[13164]=8'b11111111;
memory[13165]=8'b11111111;
memory[13166]=8'b11111111;
memory[13167]=8'b11111111;
memory[13168]=8'b11111111;
memory[13169]=8'b11111111;
memory[13170]=8'b11111111;
memory[13171]=8'b11111111;
memory[13172]=8'b11000111;
memory[13173]=8'b10000111;
memory[13174]=8'b11111111;
memory[13175]=8'b11111111;
memory[13176]=8'b11111111;
memory[13177]=8'b11111111;
memory[13178]=8'b11111111;
memory[13179]=8'b11111111;
memory[13180]=8'b11111111;
memory[13181]=8'b11111111;
memory[13182]=8'b11111111;
memory[13183]=8'b11111111;
memory[13184]=8'b11111111;
memory[13185]=8'b11111111;
memory[13186]=8'b11111111;
memory[13187]=8'b10000111;
memory[13188]=8'b10001111;
memory[13189]=8'b11111111;
memory[13190]=8'b11111111;
memory[13191]=8'b11111111;
memory[13192]=8'b11111111;
memory[13193]=8'b11111111;
memory[13194]=8'b11111111;
memory[13195]=8'b11111111;
memory[13196]=8'b11111111;
memory[13197]=8'b11111111;
memory[13198]=8'b11111111;
memory[13199]=8'b11111111;
memory[13200]=8'b11111111;
memory[13201]=8'b11111111;
memory[13202]=8'b11111111;
memory[13203]=8'b11111111;
memory[13204]=8'b11111111;
memory[13205]=8'b11111111;
memory[13206]=8'b11111111;
memory[13207]=8'b11111111;
memory[13208]=8'b11111111;
memory[13209]=8'b11111111;
memory[13210]=8'b11111111;
memory[13211]=8'b11111111;
memory[13212]=8'b11000111;
memory[13213]=8'b00001111;
memory[13214]=8'b11111111;
memory[13215]=8'b11111111;
memory[13216]=8'b11111111;
memory[13217]=8'b11111111;
memory[13218]=8'b11111111;
memory[13219]=8'b11111111;
memory[13220]=8'b11111111;
memory[13221]=8'b11111111;
memory[13222]=8'b11111111;
memory[13223]=8'b11111111;
memory[13224]=8'b11111111;
memory[13225]=8'b11111111;
memory[13226]=8'b11111111;
memory[13227]=8'b11000111;
memory[13228]=8'b10001111;
memory[13229]=8'b11111111;
memory[13230]=8'b11111111;
memory[13231]=8'b11111111;
memory[13232]=8'b11111111;
memory[13233]=8'b11111111;
memory[13234]=8'b11111111;
memory[13235]=8'b11111111;
memory[13236]=8'b11111111;
memory[13237]=8'b11111111;
memory[13238]=8'b11111111;
memory[13239]=8'b11111111;
memory[13240]=8'b11111111;
memory[13241]=8'b11111111;
memory[13242]=8'b11111111;
memory[13243]=8'b11111111;
memory[13244]=8'b11111111;
memory[13245]=8'b11111111;
memory[13246]=8'b11111111;
memory[13247]=8'b11111111;
memory[13248]=8'b11111111;
memory[13249]=8'b11111111;
memory[13250]=8'b11111111;
memory[13251]=8'b11111111;
memory[13252]=8'b11000111;
memory[13253]=8'b00001111;
memory[13254]=8'b11111111;
memory[13255]=8'b11111111;
memory[13256]=8'b11111111;
memory[13257]=8'b11111111;
memory[13258]=8'b11111111;
memory[13259]=8'b11111111;
memory[13260]=8'b11111111;
memory[13261]=8'b11111111;
memory[13262]=8'b11111111;
memory[13263]=8'b11111111;
memory[13264]=8'b11111111;
memory[13265]=8'b11111111;
memory[13266]=8'b11111111;
memory[13267]=8'b11000111;
memory[13268]=8'b10001111;
memory[13269]=8'b11111111;
memory[13270]=8'b11111111;
memory[13271]=8'b11111111;
memory[13272]=8'b11111111;
memory[13273]=8'b11111111;
memory[13274]=8'b11111111;
memory[13275]=8'b11111111;
memory[13276]=8'b11111111;
memory[13277]=8'b11111111;
memory[13278]=8'b11111111;
memory[13279]=8'b11111111;
memory[13280]=8'b11111111;
memory[13281]=8'b11111111;
memory[13282]=8'b11111111;
memory[13283]=8'b11111111;
memory[13284]=8'b11111111;
memory[13285]=8'b11111111;
memory[13286]=8'b11111111;
memory[13287]=8'b11111111;
memory[13288]=8'b11111111;
memory[13289]=8'b11111111;
memory[13290]=8'b11111111;
memory[13291]=8'b11111111;
memory[13292]=8'b10000111;
memory[13293]=8'b00001111;
memory[13294]=8'b11111111;
memory[13295]=8'b11111111;
memory[13296]=8'b11111111;
memory[13297]=8'b11111111;
memory[13298]=8'b11111111;
memory[13299]=8'b11111111;
memory[13300]=8'b11111111;
memory[13301]=8'b11111111;
memory[13302]=8'b11111111;
memory[13303]=8'b11111111;
memory[13304]=8'b11111111;
memory[13305]=8'b11111111;
memory[13306]=8'b11111111;
memory[13307]=8'b11000011;
memory[13308]=8'b10001111;
memory[13309]=8'b11111111;
memory[13310]=8'b11111111;
memory[13311]=8'b11111111;
memory[13312]=8'b11111111;
memory[13313]=8'b11111111;
memory[13314]=8'b11111111;
memory[13315]=8'b11111111;
memory[13316]=8'b11111111;
memory[13317]=8'b11111111;
memory[13318]=8'b11111111;
memory[13319]=8'b11111111;
memory[13320]=8'b11111111;
memory[13321]=8'b11111111;
memory[13322]=8'b11111111;
memory[13323]=8'b11111111;
memory[13324]=8'b11111111;
memory[13325]=8'b11111111;
memory[13326]=8'b11111111;
memory[13327]=8'b11111111;
memory[13328]=8'b11111111;
memory[13329]=8'b11111111;
memory[13330]=8'b11111111;
memory[13331]=8'b11111111;
memory[13332]=8'b10001111;
memory[13333]=8'b00000111;
memory[13334]=8'b11111111;
memory[13335]=8'b11111111;
memory[13336]=8'b11111111;
memory[13337]=8'b11111111;
memory[13338]=8'b11111111;
memory[13339]=8'b11111111;
memory[13340]=8'b11111111;
memory[13341]=8'b11111111;
memory[13342]=8'b11111111;
memory[13343]=8'b11111111;
memory[13344]=8'b11111111;
memory[13345]=8'b11111111;
memory[13346]=8'b11111111;
memory[13347]=8'b11100011;
memory[13348]=8'b11001111;
memory[13349]=8'b11111111;
memory[13350]=8'b11111111;
memory[13351]=8'b11111111;
memory[13352]=8'b11111111;
memory[13353]=8'b11111111;
memory[13354]=8'b11111111;
memory[13355]=8'b11111111;
memory[13356]=8'b11111111;
memory[13357]=8'b11111111;
memory[13358]=8'b11111111;
memory[13359]=8'b11111111;
memory[13360]=8'b11111111;
memory[13361]=8'b11111111;
memory[13362]=8'b11111111;
memory[13363]=8'b11111111;
memory[13364]=8'b11111111;
memory[13365]=8'b11111111;
memory[13366]=8'b11111111;
memory[13367]=8'b11111111;
memory[13368]=8'b11111111;
memory[13369]=8'b11111111;
memory[13370]=8'b11111111;
memory[13371]=8'b11111111;
memory[13372]=8'b10000111;
memory[13373]=8'b00000111;
memory[13374]=8'b11111111;
memory[13375]=8'b11111111;
memory[13376]=8'b11111111;
memory[13377]=8'b11111111;
memory[13378]=8'b11111111;
memory[13379]=8'b11111111;
memory[13380]=8'b11111111;
memory[13381]=8'b11111111;
memory[13382]=8'b11111111;
memory[13383]=8'b11111111;
memory[13384]=8'b11111111;
memory[13385]=8'b11111111;
memory[13386]=8'b11111111;
memory[13387]=8'b11100011;
memory[13388]=8'b11001111;
memory[13389]=8'b11111111;
memory[13390]=8'b11111111;
memory[13391]=8'b11111111;
memory[13392]=8'b11111111;
memory[13393]=8'b11111111;
memory[13394]=8'b11111111;
memory[13395]=8'b11111111;
memory[13396]=8'b11111111;
memory[13397]=8'b11111111;
memory[13398]=8'b11111111;
memory[13399]=8'b11111111;
memory[13400]=8'b11111111;
memory[13401]=8'b11111111;
memory[13402]=8'b11111111;
memory[13403]=8'b11111111;
memory[13404]=8'b11111111;
memory[13405]=8'b11111111;
memory[13406]=8'b11111111;
memory[13407]=8'b11111111;
memory[13408]=8'b11111111;
memory[13409]=8'b11111111;
memory[13410]=8'b11111111;
memory[13411]=8'b11111111;
memory[13412]=8'b10000111;
memory[13413]=8'b00000111;
memory[13414]=8'b11111111;
memory[13415]=8'b11111111;
memory[13416]=8'b11111111;
memory[13417]=8'b11111111;
memory[13418]=8'b11111111;
memory[13419]=8'b11111111;
memory[13420]=8'b11111111;
memory[13421]=8'b11111111;
memory[13422]=8'b11111111;
memory[13423]=8'b11111111;
memory[13424]=8'b11111111;
memory[13425]=8'b11111111;
memory[13426]=8'b11111111;
memory[13427]=8'b11100011;
memory[13428]=8'b11001111;
memory[13429]=8'b11111111;
memory[13430]=8'b11111111;
memory[13431]=8'b11111111;
memory[13432]=8'b11111111;
memory[13433]=8'b11111111;
memory[13434]=8'b11111111;
memory[13435]=8'b11111111;
memory[13436]=8'b11111111;
memory[13437]=8'b11111111;
memory[13438]=8'b11111111;
memory[13439]=8'b11111111;
memory[13440]=8'b11111111;
memory[13441]=8'b11111111;
memory[13442]=8'b11111111;
memory[13443]=8'b11111111;
memory[13444]=8'b11111111;
memory[13445]=8'b11111111;
memory[13446]=8'b11111111;
memory[13447]=8'b11111111;
memory[13448]=8'b11111111;
memory[13449]=8'b11111111;
memory[13450]=8'b11111111;
memory[13451]=8'b11111111;
memory[13452]=8'b00000111;
memory[13453]=8'b00000111;
memory[13454]=8'b11111111;
memory[13455]=8'b11111111;
memory[13456]=8'b11111111;
memory[13457]=8'b11111111;
memory[13458]=8'b11111111;
memory[13459]=8'b11111111;
memory[13460]=8'b11111111;
memory[13461]=8'b11111111;
memory[13462]=8'b11111111;
memory[13463]=8'b11111111;
memory[13464]=8'b11111111;
memory[13465]=8'b11111111;
memory[13466]=8'b11111111;
memory[13467]=8'b11110011;
memory[13468]=8'b11001111;
memory[13469]=8'b11111111;
memory[13470]=8'b11111111;
memory[13471]=8'b11111111;
memory[13472]=8'b11111111;
memory[13473]=8'b11111111;
memory[13474]=8'b11111111;
memory[13475]=8'b11111111;
memory[13476]=8'b11111111;
memory[13477]=8'b11111111;
memory[13478]=8'b11111111;
memory[13479]=8'b11111111;
memory[13480]=8'b11111111;
memory[13481]=8'b11111111;
memory[13482]=8'b11111111;
memory[13483]=8'b11111111;
memory[13484]=8'b11111111;
memory[13485]=8'b11111111;
memory[13486]=8'b11111111;
memory[13487]=8'b11111111;
memory[13488]=8'b11111111;
memory[13489]=8'b11111111;
memory[13490]=8'b11111111;
memory[13491]=8'b11111111;
memory[13492]=8'b00000011;
memory[13493]=8'b00000011;
memory[13494]=8'b11111111;
memory[13495]=8'b11111111;
memory[13496]=8'b11111111;
memory[13497]=8'b11111111;
memory[13498]=8'b11111111;
memory[13499]=8'b11111111;
memory[13500]=8'b11111111;
memory[13501]=8'b11111111;
memory[13502]=8'b11111111;
memory[13503]=8'b11111111;
memory[13504]=8'b11111111;
memory[13505]=8'b11111111;
memory[13506]=8'b11111111;
memory[13507]=8'b11110001;
memory[13508]=8'b11000111;
memory[13509]=8'b11111111;
memory[13510]=8'b11111111;
memory[13511]=8'b11111111;
memory[13512]=8'b11111111;
memory[13513]=8'b11111111;
memory[13514]=8'b11111111;
memory[13515]=8'b11111111;
memory[13516]=8'b11111111;
memory[13517]=8'b11111111;
memory[13518]=8'b11111111;
memory[13519]=8'b11111111;
memory[13520]=8'b11111111;
memory[13521]=8'b11111111;
memory[13522]=8'b11111111;
memory[13523]=8'b11111111;
memory[13524]=8'b11111111;
memory[13525]=8'b11111111;
memory[13526]=8'b11111111;
memory[13527]=8'b11111111;
memory[13528]=8'b11111111;
memory[13529]=8'b11111111;
memory[13530]=8'b11111111;
memory[13531]=8'b11111111;
memory[13532]=8'b00000001;
memory[13533]=8'b00000011;
memory[13534]=8'b11111111;
memory[13535]=8'b11111111;
memory[13536]=8'b11111111;
memory[13537]=8'b11111111;
memory[13538]=8'b11111111;
memory[13539]=8'b11111111;
memory[13540]=8'b11111111;
memory[13541]=8'b11111111;
memory[13542]=8'b11111111;
memory[13543]=8'b11111111;
memory[13544]=8'b11111111;
memory[13545]=8'b11111111;
memory[13546]=8'b11111111;
memory[13547]=8'b11110001;
memory[13548]=8'b11100111;
memory[13549]=8'b11111111;
memory[13550]=8'b11111111;
memory[13551]=8'b11111111;
memory[13552]=8'b11111111;
memory[13553]=8'b11111111;
memory[13554]=8'b11111111;
memory[13555]=8'b11111111;
memory[13556]=8'b11111111;
memory[13557]=8'b11111111;
memory[13558]=8'b11111111;
memory[13559]=8'b11111111;
memory[13560]=8'b11111111;
memory[13561]=8'b11111111;
memory[13562]=8'b11111111;
memory[13563]=8'b11111111;
memory[13564]=8'b11111111;
memory[13565]=8'b11111111;
memory[13566]=8'b11111111;
memory[13567]=8'b11111111;
memory[13568]=8'b11111111;
memory[13569]=8'b11111111;
memory[13570]=8'b11111111;
memory[13571]=8'b11111111;
memory[13572]=8'b10000001;
memory[13573]=8'b10000111;
memory[13574]=8'b11111111;
memory[13575]=8'b11111111;
memory[13576]=8'b11111111;
memory[13577]=8'b11111111;
memory[13578]=8'b11111111;
memory[13579]=8'b11111111;
memory[13580]=8'b11111111;
memory[13581]=8'b11111111;
memory[13582]=8'b11111111;
memory[13583]=8'b11111111;
memory[13584]=8'b11111111;
memory[13585]=8'b11111111;
memory[13586]=8'b11111111;
memory[13587]=8'b11110001;
memory[13588]=8'b11100111;
memory[13589]=8'b11111111;
memory[13590]=8'b11111111;
memory[13591]=8'b11111111;
memory[13592]=8'b11111111;
memory[13593]=8'b11111111;
memory[13594]=8'b11111111;
memory[13595]=8'b11111111;
memory[13596]=8'b11111111;
memory[13597]=8'b11111111;
memory[13598]=8'b11111111;
memory[13599]=8'b11111111;
memory[13600]=8'b11111111;
memory[13601]=8'b11111111;
memory[13602]=8'b11111111;
memory[13603]=8'b11111111;
memory[13604]=8'b11111111;
memory[13605]=8'b11111111;
memory[13606]=8'b11111111;
memory[13607]=8'b11111111;
memory[13608]=8'b11111111;
memory[13609]=8'b11111111;
memory[13610]=8'b11111111;
memory[13611]=8'b11111111;
memory[13612]=8'b10000001;
memory[13613]=8'b10000111;
memory[13614]=8'b11111111;
memory[13615]=8'b11111111;
memory[13616]=8'b11111111;
memory[13617]=8'b11111111;
memory[13618]=8'b11111111;
memory[13619]=8'b11111111;
memory[13620]=8'b11111111;
memory[13621]=8'b11111111;
memory[13622]=8'b11111111;
memory[13623]=8'b11111111;
memory[13624]=8'b11111111;
memory[13625]=8'b11111111;
memory[13626]=8'b11111111;
memory[13627]=8'b11110001;
memory[13628]=8'b11100111;
memory[13629]=8'b11111111;
memory[13630]=8'b11111111;
memory[13631]=8'b11111111;
memory[13632]=8'b11111111;
memory[13633]=8'b11111111;
memory[13634]=8'b11111111;
memory[13635]=8'b11111111;
memory[13636]=8'b11111111;
memory[13637]=8'b11111111;
memory[13638]=8'b11111111;
memory[13639]=8'b11111111;
memory[13640]=8'b11111111;
memory[13641]=8'b11111111;
memory[13642]=8'b11111111;
memory[13643]=8'b11111111;
memory[13644]=8'b11111111;
memory[13645]=8'b11111111;
memory[13646]=8'b11111111;
memory[13647]=8'b11111111;
memory[13648]=8'b11111111;
memory[13649]=8'b11111111;
memory[13650]=8'b11111111;
memory[13651]=8'b11111111;
memory[13652]=8'b11000001;
memory[13653]=8'b10000111;
memory[13654]=8'b11111111;
memory[13655]=8'b11111111;
memory[13656]=8'b11111111;
memory[13657]=8'b11111111;
memory[13658]=8'b11111111;
memory[13659]=8'b11111111;
memory[13660]=8'b11111111;
memory[13661]=8'b11111111;
memory[13662]=8'b11111111;
memory[13663]=8'b11111111;
memory[13664]=8'b11111111;
memory[13665]=8'b11111111;
memory[13666]=8'b11111111;
memory[13667]=8'b11111000;
memory[13668]=8'b11100111;
memory[13669]=8'b11111111;
memory[13670]=8'b11111111;
memory[13671]=8'b11111111;
memory[13672]=8'b11111111;
memory[13673]=8'b11111111;
memory[13674]=8'b11111111;
memory[13675]=8'b11111111;
memory[13676]=8'b11111111;
memory[13677]=8'b11111111;
memory[13678]=8'b11111111;
memory[13679]=8'b11111111;
memory[13680]=8'b11111111;
memory[13681]=8'b11111111;
memory[13682]=8'b11111111;
memory[13683]=8'b11111111;
memory[13684]=8'b11111111;
memory[13685]=8'b11111111;
memory[13686]=8'b11111111;
memory[13687]=8'b11111111;
memory[13688]=8'b11111111;
memory[13689]=8'b11111111;
memory[13690]=8'b11111111;
memory[13691]=8'b11111111;
memory[13692]=8'b11100001;
memory[13693]=8'b10000111;
memory[13694]=8'b11111111;
memory[13695]=8'b11111111;
memory[13696]=8'b11111111;
memory[13697]=8'b11111111;
memory[13698]=8'b11111111;
memory[13699]=8'b11111111;
memory[13700]=8'b11111111;
memory[13701]=8'b11111111;
memory[13702]=8'b11111111;
memory[13703]=8'b11111111;
memory[13704]=8'b11111111;
memory[13705]=8'b11111111;
memory[13706]=8'b11111111;
memory[13707]=8'b11111000;
memory[13708]=8'b11100111;
memory[13709]=8'b11111111;
memory[13710]=8'b11111111;
memory[13711]=8'b11111111;
memory[13712]=8'b11111111;
memory[13713]=8'b11111111;
memory[13714]=8'b11111111;
memory[13715]=8'b11111111;
memory[13716]=8'b11111111;
memory[13717]=8'b11111111;
memory[13718]=8'b11111111;
memory[13719]=8'b11111111;
memory[13720]=8'b11111111;
memory[13721]=8'b11111111;
memory[13722]=8'b11111111;
memory[13723]=8'b11111111;
memory[13724]=8'b11111111;
memory[13725]=8'b11111111;
memory[13726]=8'b11111111;
memory[13727]=8'b11111111;
memory[13728]=8'b11111111;
memory[13729]=8'b11111111;
memory[13730]=8'b11111111;
memory[13731]=8'b11111111;
memory[13732]=8'b11100001;
memory[13733]=8'b10000111;
memory[13734]=8'b11111111;
memory[13735]=8'b11111111;
memory[13736]=8'b11111111;
memory[13737]=8'b11111111;
memory[13738]=8'b11111111;
memory[13739]=8'b11111111;
memory[13740]=8'b11111111;
memory[13741]=8'b11111111;
memory[13742]=8'b11111111;
memory[13743]=8'b11111111;
memory[13744]=8'b11111111;
memory[13745]=8'b11111111;
memory[13746]=8'b11111111;
memory[13747]=8'b11111000;
memory[13748]=8'b11100111;
memory[13749]=8'b11111111;
memory[13750]=8'b11111111;
memory[13751]=8'b11111111;
memory[13752]=8'b11111111;
memory[13753]=8'b11111111;
memory[13754]=8'b11111111;
memory[13755]=8'b11111111;
memory[13756]=8'b11111111;
memory[13757]=8'b11111111;
memory[13758]=8'b11111111;
memory[13759]=8'b11111111;
memory[13760]=8'b11111111;
memory[13761]=8'b11111111;
memory[13762]=8'b11111111;
memory[13763]=8'b11111111;
memory[13764]=8'b11111111;
memory[13765]=8'b11111111;
memory[13766]=8'b11111111;
memory[13767]=8'b11111111;
memory[13768]=8'b11111111;
memory[13769]=8'b11111111;
memory[13770]=8'b11111111;
memory[13771]=8'b11111111;
memory[13772]=8'b11110000;
memory[13773]=8'b11000111;
memory[13774]=8'b11111111;
memory[13775]=8'b11111111;
memory[13776]=8'b11111111;
memory[13777]=8'b11111111;
memory[13778]=8'b11111111;
memory[13779]=8'b11111111;
memory[13780]=8'b11111111;
memory[13781]=8'b11111111;
memory[13782]=8'b11111111;
memory[13783]=8'b11111111;
memory[13784]=8'b11111111;
memory[13785]=8'b11111111;
memory[13786]=8'b11111111;
memory[13787]=8'b11111100;
memory[13788]=8'b01110011;
memory[13789]=8'b11111111;
memory[13790]=8'b11111111;
memory[13791]=8'b11111111;
memory[13792]=8'b11111111;
memory[13793]=8'b11111111;
memory[13794]=8'b11111111;
memory[13795]=8'b11111111;
memory[13796]=8'b11111111;
memory[13797]=8'b11111111;
memory[13798]=8'b11111111;
memory[13799]=8'b11111111;
memory[13800]=8'b11111111;
memory[13801]=8'b11111111;
memory[13802]=8'b11111111;
memory[13803]=8'b11111111;
memory[13804]=8'b11111111;
memory[13805]=8'b11111111;
memory[13806]=8'b11111111;
memory[13807]=8'b11111111;
memory[13808]=8'b11111111;
memory[13809]=8'b11111111;
memory[13810]=8'b11111111;
memory[13811]=8'b11111111;
memory[13812]=8'b11110000;
memory[13813]=8'b11000111;
memory[13814]=8'b11111111;
memory[13815]=8'b11111111;
memory[13816]=8'b11111111;
memory[13817]=8'b11111111;
memory[13818]=8'b11111111;
memory[13819]=8'b11111111;
memory[13820]=8'b11111111;
memory[13821]=8'b11111111;
memory[13822]=8'b11111111;
memory[13823]=8'b11111111;
memory[13824]=8'b11111111;
memory[13825]=8'b11111111;
memory[13826]=8'b11111111;
memory[13827]=8'b11111100;
memory[13828]=8'b01110011;
memory[13829]=8'b11111111;
memory[13830]=8'b11111111;
memory[13831]=8'b11111111;
memory[13832]=8'b11111111;
memory[13833]=8'b11111111;
memory[13834]=8'b11111111;
memory[13835]=8'b11111111;
memory[13836]=8'b11111111;
memory[13837]=8'b11111111;
memory[13838]=8'b11111111;
memory[13839]=8'b11111111;
memory[13840]=8'b11111111;
memory[13841]=8'b11111111;
memory[13842]=8'b11111111;
memory[13843]=8'b11111111;
memory[13844]=8'b11111111;
memory[13845]=8'b11111111;
memory[13846]=8'b11111111;
memory[13847]=8'b11111111;
memory[13848]=8'b11111111;
memory[13849]=8'b11111111;
memory[13850]=8'b11111111;
memory[13851]=8'b11111111;
memory[13852]=8'b11111000;
memory[13853]=8'b11100111;
memory[13854]=8'b11111111;
memory[13855]=8'b11111111;
memory[13856]=8'b11111111;
memory[13857]=8'b11111111;
memory[13858]=8'b11111111;
memory[13859]=8'b11111111;
memory[13860]=8'b11111111;
memory[13861]=8'b11111111;
memory[13862]=8'b11111111;
memory[13863]=8'b11111111;
memory[13864]=8'b11110011;
memory[13865]=8'b11111111;
memory[13866]=8'b11111111;
memory[13867]=8'b11111100;
memory[13868]=8'b01110011;
memory[13869]=8'b11111111;
memory[13870]=8'b11111111;
memory[13871]=8'b11111111;
memory[13872]=8'b11111111;
memory[13873]=8'b11111111;
memory[13874]=8'b11111111;
memory[13875]=8'b11111111;
memory[13876]=8'b11111111;
memory[13877]=8'b11111111;
memory[13878]=8'b11111111;
memory[13879]=8'b11111111;
memory[13880]=8'b11111111;
memory[13881]=8'b11111111;
memory[13882]=8'b11111111;
memory[13883]=8'b11111111;
memory[13884]=8'b11111111;
memory[13885]=8'b11111111;
memory[13886]=8'b11111111;
memory[13887]=8'b11111111;
memory[13888]=8'b11111111;
memory[13889]=8'b11111111;
memory[13890]=8'b11111111;
memory[13891]=8'b11111111;
memory[13892]=8'b11111000;
memory[13893]=8'b01100111;
memory[13894]=8'b11111111;
memory[13895]=8'b11111111;
memory[13896]=8'b11111111;
memory[13897]=8'b11111111;
memory[13898]=8'b11111111;
memory[13899]=8'b11111111;
memory[13900]=8'b11111111;
memory[13901]=8'b11111111;
memory[13902]=8'b11111111;
memory[13903]=8'b11111111;
memory[13904]=8'b11100000;
memory[13905]=8'b01111111;
memory[13906]=8'b11111111;
memory[13907]=8'b11111100;
memory[13908]=8'b01110011;
memory[13909]=8'b11111111;
memory[13910]=8'b11111111;
memory[13911]=8'b11111111;
memory[13912]=8'b11111111;
memory[13913]=8'b11111111;
memory[13914]=8'b11111111;
memory[13915]=8'b11111111;
memory[13916]=8'b11111111;
memory[13917]=8'b11111111;
memory[13918]=8'b11111111;
memory[13919]=8'b11111111;
memory[13920]=8'b11111111;
memory[13921]=8'b11111111;
memory[13922]=8'b11111111;
memory[13923]=8'b11111111;
memory[13924]=8'b11111111;
memory[13925]=8'b11111111;
memory[13926]=8'b11111111;
memory[13927]=8'b11111111;
memory[13928]=8'b11111111;
memory[13929]=8'b11111111;
memory[13930]=8'b11111111;
memory[13931]=8'b11111111;
memory[13932]=8'b11111100;
memory[13933]=8'b01111111;
memory[13934]=8'b11111111;
memory[13935]=8'b11111111;
memory[13936]=8'b11111111;
memory[13937]=8'b11111111;
memory[13938]=8'b11111111;
memory[13939]=8'b11111111;
memory[13940]=8'b11111111;
memory[13941]=8'b11111111;
memory[13942]=8'b11111111;
memory[13943]=8'b11111111;
memory[13944]=8'b11000011;
memory[13945]=8'b11111111;
memory[13946]=8'b11111111;
memory[13947]=8'b11111100;
memory[13948]=8'b01110001;
memory[13949]=8'b11111111;
memory[13950]=8'b11111111;
memory[13951]=8'b11111111;
memory[13952]=8'b11111111;
memory[13953]=8'b11111111;
memory[13954]=8'b11111111;
memory[13955]=8'b11111111;
memory[13956]=8'b11111111;
memory[13957]=8'b11111111;
memory[13958]=8'b11111111;
memory[13959]=8'b11111111;
memory[13960]=8'b11111111;
memory[13961]=8'b11111111;
memory[13962]=8'b11111111;
memory[13963]=8'b11111111;
memory[13964]=8'b11111111;
memory[13965]=8'b11111111;
memory[13966]=8'b11111111;
memory[13967]=8'b11111111;
memory[13968]=8'b11111111;
memory[13969]=8'b11111111;
memory[13970]=8'b11111111;
memory[13971]=8'b11111111;
memory[13972]=8'b11111100;
memory[13973]=8'b00111111;
memory[13974]=8'b11111111;
memory[13975]=8'b11111111;
memory[13976]=8'b11111111;
memory[13977]=8'b11111111;
memory[13978]=8'b11111111;
memory[13979]=8'b11111111;
memory[13980]=8'b11111111;
memory[13981]=8'b11111111;
memory[13982]=8'b11111111;
memory[13983]=8'b11111111;
memory[13984]=8'b11001111;
memory[13985]=8'b11111111;
memory[13986]=8'b11111111;
memory[13987]=8'b11111100;
memory[13988]=8'b01110001;
memory[13989]=8'b11111111;
memory[13990]=8'b11111111;
memory[13991]=8'b11111111;
memory[13992]=8'b11111111;
memory[13993]=8'b11111111;
memory[13994]=8'b11111111;
memory[13995]=8'b11111111;
memory[13996]=8'b11111111;
memory[13997]=8'b11111111;
memory[13998]=8'b11111111;
memory[13999]=8'b11111111;
memory[14000]=8'b11111111;
memory[14001]=8'b11111111;
memory[14002]=8'b11111111;
memory[14003]=8'b11111111;
memory[14004]=8'b11111111;
memory[14005]=8'b11111111;
memory[14006]=8'b11111111;
memory[14007]=8'b11111111;
memory[14008]=8'b11111111;
memory[14009]=8'b11111111;
memory[14010]=8'b11111111;
memory[14011]=8'b11111111;
memory[14012]=8'b11111110;
memory[14013]=8'b00011111;
memory[14014]=8'b11111111;
memory[14015]=8'b11111111;
memory[14016]=8'b11111111;
memory[14017]=8'b11111111;
memory[14018]=8'b11111111;
memory[14019]=8'b11111111;
memory[14020]=8'b11111111;
memory[14021]=8'b11111111;
memory[14022]=8'b11111111;
memory[14023]=8'b11111111;
memory[14024]=8'b10011111;
memory[14025]=8'b11111111;
memory[14026]=8'b11111111;
memory[14027]=8'b11111000;
memory[14028]=8'b01100001;
memory[14029]=8'b11111111;
memory[14030]=8'b11111111;
memory[14031]=8'b11111111;
memory[14032]=8'b11111111;
memory[14033]=8'b11111111;
memory[14034]=8'b11111111;
memory[14035]=8'b11111111;
memory[14036]=8'b11111111;
memory[14037]=8'b11111111;
memory[14038]=8'b11111111;
memory[14039]=8'b11111111;
memory[14040]=8'b11111111;
memory[14041]=8'b11111111;
memory[14042]=8'b11111111;
memory[14043]=8'b11111111;
memory[14044]=8'b11111111;
memory[14045]=8'b11111111;
memory[14046]=8'b11111111;
memory[14047]=8'b11111111;
memory[14048]=8'b11111111;
memory[14049]=8'b11111111;
memory[14050]=8'b11111111;
memory[14051]=8'b11111111;
memory[14052]=8'b11111110;
memory[14053]=8'b00011111;
memory[14054]=8'b11111111;
memory[14055]=8'b11111111;
memory[14056]=8'b11111111;
memory[14057]=8'b11111111;
memory[14058]=8'b11111111;
memory[14059]=8'b11111111;
memory[14060]=8'b11111111;
memory[14061]=8'b11111111;
memory[14062]=8'b10000111;
memory[14063]=8'b11111111;
memory[14064]=8'b10111111;
memory[14065]=8'b11111111;
memory[14066]=8'b11111111;
memory[14067]=8'b11111000;
memory[14068]=8'b01100000;
memory[14069]=8'b11111111;
memory[14070]=8'b11111111;
memory[14071]=8'b11111111;
memory[14072]=8'b11111111;
memory[14073]=8'b11111111;
memory[14074]=8'b11111111;
memory[14075]=8'b11111111;
memory[14076]=8'b11111111;
memory[14077]=8'b11111111;
memory[14078]=8'b11111111;
memory[14079]=8'b11111111;
memory[14080]=8'b11111111;
memory[14081]=8'b11111111;
memory[14082]=8'b11111111;
memory[14083]=8'b11111111;
memory[14084]=8'b11111111;
memory[14085]=8'b11111111;
memory[14086]=8'b11111111;
memory[14087]=8'b11111111;
memory[14088]=8'b11111111;
memory[14089]=8'b11111111;
memory[14090]=8'b11111111;
memory[14091]=8'b11111111;
memory[14092]=8'b11111111;
memory[14093]=8'b00011111;
memory[14094]=8'b11111111;
memory[14095]=8'b11111111;
memory[14096]=8'b11111111;
memory[14097]=8'b11111111;
memory[14098]=8'b11111111;
memory[14099]=8'b11111111;
memory[14100]=8'b11111111;
memory[14101]=8'b11111111;
memory[14102]=8'b11111111;
memory[14103]=8'b11111111;
memory[14104]=8'b11111111;
memory[14105]=8'b11111111;
memory[14106]=8'b11111111;
memory[14107]=8'b11111000;
memory[14108]=8'b01100001;
memory[14109]=8'b11111111;
memory[14110]=8'b11111111;
memory[14111]=8'b11111111;
memory[14112]=8'b11111111;
memory[14113]=8'b11111111;
memory[14114]=8'b11111111;
memory[14115]=8'b11111111;
memory[14116]=8'b11111111;
memory[14117]=8'b11111111;
memory[14118]=8'b11111111;
memory[14119]=8'b11111111;
memory[14120]=8'b11111111;
memory[14121]=8'b11111111;
memory[14122]=8'b11111111;
memory[14123]=8'b11111111;
memory[14124]=8'b11111111;
memory[14125]=8'b11111111;
memory[14126]=8'b11111111;
memory[14127]=8'b11111111;
memory[14128]=8'b11111111;
memory[14129]=8'b11111111;
memory[14130]=8'b11111111;
memory[14131]=8'b11111111;
memory[14132]=8'b11111111;
memory[14133]=8'b00001111;
memory[14134]=8'b11111111;
memory[14135]=8'b11111111;
memory[14136]=8'b11111111;
memory[14137]=8'b11111111;
memory[14138]=8'b11111111;
memory[14139]=8'b11111111;
memory[14140]=8'b11111111;
memory[14141]=8'b11111111;
memory[14142]=8'b11111111;
memory[14143]=8'b11111111;
memory[14144]=8'b11111111;
memory[14145]=8'b11111111;
memory[14146]=8'b11111111;
memory[14147]=8'b11111000;
memory[14148]=8'b01000001;
memory[14149]=8'b11111111;
memory[14150]=8'b11111111;
memory[14151]=8'b11111111;
memory[14152]=8'b11111111;
memory[14153]=8'b11111111;
memory[14154]=8'b11111111;
memory[14155]=8'b11111111;
memory[14156]=8'b11111111;
memory[14157]=8'b11111111;
memory[14158]=8'b11111111;
memory[14159]=8'b11111111;
memory[14160]=8'b11111111;
memory[14161]=8'b11111111;
memory[14162]=8'b11111111;
memory[14163]=8'b11111111;
memory[14164]=8'b11111111;
memory[14165]=8'b11111111;
memory[14166]=8'b11111111;
memory[14167]=8'b11111111;
memory[14168]=8'b11111111;
memory[14169]=8'b11111111;
memory[14170]=8'b11111111;
memory[14171]=8'b11111111;
memory[14172]=8'b11111111;
memory[14173]=8'b10001111;
memory[14174]=8'b11111111;
memory[14175]=8'b11111111;
memory[14176]=8'b11111111;
memory[14177]=8'b11111111;
memory[14178]=8'b11111111;
memory[14179]=8'b11111111;
memory[14180]=8'b11111111;
memory[14181]=8'b11111111;
memory[14182]=8'b11111101;
memory[14183]=8'b11111111;
memory[14184]=8'b11111111;
memory[14185]=8'b11111111;
memory[14186]=8'b11111111;
memory[14187]=8'b11111100;
memory[14188]=8'b01000011;
memory[14189]=8'b11111111;
memory[14190]=8'b11111111;
memory[14191]=8'b11111111;
memory[14192]=8'b11111111;
memory[14193]=8'b11111111;
memory[14194]=8'b11111111;
memory[14195]=8'b11111111;
memory[14196]=8'b11111111;
memory[14197]=8'b11111111;
memory[14198]=8'b11111111;
memory[14199]=8'b11111111;
memory[14200]=8'b11111111;
memory[14201]=8'b11111111;
memory[14202]=8'b11111111;
memory[14203]=8'b11111111;
memory[14204]=8'b11111111;
memory[14205]=8'b11111111;
memory[14206]=8'b11111111;
memory[14207]=8'b11111111;
memory[14208]=8'b11111111;
memory[14209]=8'b11111111;
memory[14210]=8'b11111111;
memory[14211]=8'b11111111;
memory[14212]=8'b11111111;
memory[14213]=8'b10001111;
memory[14214]=8'b11111111;
memory[14215]=8'b11111111;
memory[14216]=8'b11111111;
memory[14217]=8'b11111111;
memory[14218]=8'b11111111;
memory[14219]=8'b11111111;
memory[14220]=8'b11111111;
memory[14221]=8'b11111111;
memory[14222]=8'b11111000;
memory[14223]=8'b00111111;
memory[14224]=8'b11111001;
memory[14225]=8'b11111111;
memory[14226]=8'b11111111;
memory[14227]=8'b11111100;
memory[14228]=8'b10000111;
memory[14229]=8'b11111111;
memory[14230]=8'b11111111;
memory[14231]=8'b11111111;
memory[14232]=8'b11111111;
memory[14233]=8'b11111111;
memory[14234]=8'b11111111;
memory[14235]=8'b11111111;
memory[14236]=8'b11111111;
memory[14237]=8'b11111111;
memory[14238]=8'b11111111;
memory[14239]=8'b11111111;
memory[14240]=8'b11111111;
memory[14241]=8'b11111111;
memory[14242]=8'b11111111;
memory[14243]=8'b11111111;
memory[14244]=8'b11111111;
memory[14245]=8'b11111111;
memory[14246]=8'b11111111;
memory[14247]=8'b11111111;
memory[14248]=8'b11111111;
memory[14249]=8'b11111111;
memory[14250]=8'b11111111;
memory[14251]=8'b11111111;
memory[14252]=8'b11111111;
memory[14253]=8'b11000111;
memory[14254]=8'b11111111;
memory[14255]=8'b11111111;
memory[14256]=8'b11111111;
memory[14257]=8'b11111111;
memory[14258]=8'b11111111;
memory[14259]=8'b11111111;
memory[14260]=8'b11111111;
memory[14261]=8'b11111111;
memory[14262]=8'b11111110;
memory[14263]=8'b00001111;
memory[14264]=8'b11111011;
memory[14265]=8'b11111111;
memory[14266]=8'b11111111;
memory[14267]=8'b11111100;
memory[14268]=8'b10000111;
memory[14269]=8'b11111111;
memory[14270]=8'b11111111;
memory[14271]=8'b11111111;
memory[14272]=8'b11111111;
memory[14273]=8'b11111111;
memory[14274]=8'b11111111;
memory[14275]=8'b11111111;
memory[14276]=8'b11111111;
memory[14277]=8'b11111111;
memory[14278]=8'b11111111;
memory[14279]=8'b11111111;
memory[14280]=8'b11111111;
memory[14281]=8'b11111111;
memory[14282]=8'b11111111;
memory[14283]=8'b11111111;
memory[14284]=8'b11111111;
memory[14285]=8'b11111111;
memory[14286]=8'b11111111;
memory[14287]=8'b11111111;
memory[14288]=8'b11111111;
memory[14289]=8'b11111111;
memory[14290]=8'b11111111;
memory[14291]=8'b11111111;
memory[14292]=8'b11111111;
memory[14293]=8'b11000111;
memory[14294]=8'b11111111;
memory[14295]=8'b11111111;
memory[14296]=8'b11111111;
memory[14297]=8'b11111111;
memory[14298]=8'b11111111;
memory[14299]=8'b11111111;
memory[14300]=8'b11111111;
memory[14301]=8'b11111111;
memory[14302]=8'b11111111;
memory[14303]=8'b10000111;
memory[14304]=8'b11111111;
memory[14305]=8'b11111111;
memory[14306]=8'b11111111;
memory[14307]=8'b11111100;
memory[14308]=8'b10001111;
memory[14309]=8'b11111111;
memory[14310]=8'b11111111;
memory[14311]=8'b11111111;
memory[14312]=8'b11111111;
memory[14313]=8'b11111111;
memory[14314]=8'b11111111;
memory[14315]=8'b11111111;
memory[14316]=8'b11111111;
memory[14317]=8'b11111111;
memory[14318]=8'b11111111;
memory[14319]=8'b11111111;
memory[14320]=8'b11111111;
memory[14321]=8'b11111111;
memory[14322]=8'b11111111;
memory[14323]=8'b11111111;
memory[14324]=8'b11111111;
memory[14325]=8'b11111111;
memory[14326]=8'b11111111;
memory[14327]=8'b11111111;
memory[14328]=8'b11111111;
memory[14329]=8'b11111111;
memory[14330]=8'b11111111;
memory[14331]=8'b11111111;
memory[14332]=8'b11111111;
memory[14333]=8'b11000111;
memory[14334]=8'b11111111;
memory[14335]=8'b11111111;
memory[14336]=8'b11111111;
memory[14337]=8'b11111111;
memory[14338]=8'b11111111;
memory[14339]=8'b11111111;
memory[14340]=8'b11111111;
memory[14341]=8'b11111111;
memory[14342]=8'b11111110;
memory[14343]=8'b00000001;
memory[14344]=8'b11111111;
memory[14345]=8'b11111111;
memory[14346]=8'b11111111;
memory[14347]=8'b11111000;
memory[14348]=8'b00001111;
memory[14349]=8'b11111111;
memory[14350]=8'b11111111;
memory[14351]=8'b11111111;
memory[14352]=8'b11111111;
memory[14353]=8'b11111111;
memory[14354]=8'b11111111;
memory[14355]=8'b11111111;
memory[14356]=8'b11111111;
memory[14357]=8'b11111111;
memory[14358]=8'b11111111;
memory[14359]=8'b11111111;
memory[14360]=8'b11111111;
memory[14361]=8'b11111111;
memory[14362]=8'b11111111;
memory[14363]=8'b11111111;
memory[14364]=8'b11111111;
memory[14365]=8'b11111111;
memory[14366]=8'b11111111;
memory[14367]=8'b11111111;
memory[14368]=8'b11111111;
memory[14369]=8'b11111111;
memory[14370]=8'b11111111;
memory[14371]=8'b11111111;
memory[14372]=8'b11111111;
memory[14373]=8'b11100011;
memory[14374]=8'b11111111;
memory[14375]=8'b11111111;
memory[14376]=8'b11111111;
memory[14377]=8'b11111111;
memory[14378]=8'b11111111;
memory[14379]=8'b11111111;
memory[14380]=8'b11111111;
memory[14381]=8'b11111111;
memory[14382]=8'b11111111;
memory[14383]=8'b10000000;
memory[14384]=8'b11111111;
memory[14385]=8'b11111111;
memory[14386]=8'b11111111;
memory[14387]=8'b11111111;
memory[14388]=8'b00011111;
memory[14389]=8'b11111111;
memory[14390]=8'b11111111;
memory[14391]=8'b11111111;
memory[14392]=8'b11111111;
memory[14393]=8'b11111111;
memory[14394]=8'b11111111;
memory[14395]=8'b11111111;
memory[14396]=8'b11111111;
memory[14397]=8'b11111111;
memory[14398]=8'b11111111;
memory[14399]=8'b11111111;
memory[14400]=8'b11111111;
memory[14401]=8'b11111111;
memory[14402]=8'b11111111;
memory[14403]=8'b11111111;
memory[14404]=8'b11111111;
memory[14405]=8'b11111111;
memory[14406]=8'b11111111;
memory[14407]=8'b11111111;
memory[14408]=8'b11111111;
memory[14409]=8'b11111111;
memory[14410]=8'b11111111;
memory[14411]=8'b11111111;
memory[14412]=8'b11111111;
memory[14413]=8'b11100011;
memory[14414]=8'b11111111;
memory[14415]=8'b11111111;
memory[14416]=8'b11111111;
memory[14417]=8'b11111111;
memory[14418]=8'b11111111;
memory[14419]=8'b11111111;
memory[14420]=8'b11111111;
memory[14421]=8'b11111111;
memory[14422]=8'b11111111;
memory[14423]=8'b11111000;
memory[14424]=8'b11111111;
memory[14425]=8'b11111111;
memory[14426]=8'b11111111;
memory[14427]=8'b11111111;
memory[14428]=8'b00011111;
memory[14429]=8'b11111111;
memory[14430]=8'b11111111;
memory[14431]=8'b11111111;
memory[14432]=8'b11111111;
memory[14433]=8'b11111111;
memory[14434]=8'b11111111;
memory[14435]=8'b11111111;
memory[14436]=8'b11111111;
memory[14437]=8'b11111111;
memory[14438]=8'b11111111;
memory[14439]=8'b11111111;
memory[14440]=8'b11111111;
memory[14441]=8'b11111111;
memory[14442]=8'b11111111;
memory[14443]=8'b11111111;
memory[14444]=8'b11111111;
memory[14445]=8'b11111111;
memory[14446]=8'b11111111;
memory[14447]=8'b11111111;
memory[14448]=8'b11111111;
memory[14449]=8'b11111111;
memory[14450]=8'b11111111;
memory[14451]=8'b11111111;
memory[14452]=8'b11111111;
memory[14453]=8'b11110011;
memory[14454]=8'b11111111;
memory[14455]=8'b11111111;
memory[14456]=8'b11111111;
memory[14457]=8'b11111111;
memory[14458]=8'b11111111;
memory[14459]=8'b11111111;
memory[14460]=8'b11111111;
memory[14461]=8'b11111111;
memory[14462]=8'b11111111;
memory[14463]=8'b11111110;
memory[14464]=8'b01111111;
memory[14465]=8'b11111111;
memory[14466]=8'b11111111;
memory[14467]=8'b11111110;
memory[14468]=8'b00111111;
memory[14469]=8'b11111111;
memory[14470]=8'b11111111;
memory[14471]=8'b11111111;
memory[14472]=8'b11111111;
memory[14473]=8'b11111111;
memory[14474]=8'b11111111;
memory[14475]=8'b11111111;
memory[14476]=8'b11111111;
memory[14477]=8'b11111111;
memory[14478]=8'b11111111;
memory[14479]=8'b11111111;
memory[14480]=8'b11111111;
memory[14481]=8'b11111111;
memory[14482]=8'b11111111;
memory[14483]=8'b11111111;
memory[14484]=8'b11111111;
memory[14485]=8'b11111111;
memory[14486]=8'b11111111;
memory[14487]=8'b11111111;
memory[14488]=8'b11111111;
memory[14489]=8'b11111111;
memory[14490]=8'b11111111;
memory[14491]=8'b11111111;
memory[14492]=8'b11111111;
memory[14493]=8'b11110011;
memory[14494]=8'b11111111;
memory[14495]=8'b11111111;
memory[14496]=8'b11111111;
memory[14497]=8'b11111111;
memory[14498]=8'b11111111;
memory[14499]=8'b11111111;
memory[14500]=8'b11111111;
memory[14501]=8'b11111111;
memory[14502]=8'b11111111;
memory[14503]=8'b11111111;
memory[14504]=8'b00111111;
memory[14505]=8'b11111111;
memory[14506]=8'b11111111;
memory[14507]=8'b11111110;
memory[14508]=8'b00111111;
memory[14509]=8'b11111111;
memory[14510]=8'b11111111;
memory[14511]=8'b11111111;
memory[14512]=8'b11111111;
memory[14513]=8'b11111111;
memory[14514]=8'b11111111;
memory[14515]=8'b11111111;
memory[14516]=8'b11111111;
memory[14517]=8'b11111111;
memory[14518]=8'b11111111;
memory[14519]=8'b11111111;
memory[14520]=8'b11111111;
memory[14521]=8'b11111111;
memory[14522]=8'b11111111;
memory[14523]=8'b11111111;
memory[14524]=8'b11111111;
memory[14525]=8'b11111111;
memory[14526]=8'b11111111;
memory[14527]=8'b11111111;
memory[14528]=8'b11111111;
memory[14529]=8'b11111111;
memory[14530]=8'b11111111;
memory[14531]=8'b11111111;
memory[14532]=8'b11111111;
memory[14533]=8'b11110001;
memory[14534]=8'b11111111;
memory[14535]=8'b11111111;
memory[14536]=8'b11111111;
memory[14537]=8'b11111111;
memory[14538]=8'b11111111;
memory[14539]=8'b11111111;
memory[14540]=8'b11111111;
memory[14541]=8'b11111111;
memory[14542]=8'b11111111;
memory[14543]=8'b11111111;
memory[14544]=8'b00111111;
memory[14545]=8'b11111111;
memory[14546]=8'b11111111;
memory[14547]=8'b11111110;
memory[14548]=8'b01111111;
memory[14549]=8'b11111111;
memory[14550]=8'b11111111;
memory[14551]=8'b11111111;
memory[14552]=8'b11111111;
memory[14553]=8'b11111111;
memory[14554]=8'b11111111;
memory[14555]=8'b11111111;
memory[14556]=8'b11111111;
memory[14557]=8'b11111111;
memory[14558]=8'b11111111;
memory[14559]=8'b11111111;
memory[14560]=8'b11111111;
memory[14561]=8'b11111111;
memory[14562]=8'b11111111;
memory[14563]=8'b11111111;
memory[14564]=8'b11111111;
memory[14565]=8'b11111111;
memory[14566]=8'b11111111;
memory[14567]=8'b11111111;
memory[14568]=8'b11111111;
memory[14569]=8'b11111111;
memory[14570]=8'b11111111;
memory[14571]=8'b11111111;
memory[14572]=8'b11111111;
memory[14573]=8'b11111001;
memory[14574]=8'b11111111;
memory[14575]=8'b11111111;
memory[14576]=8'b11111111;
memory[14577]=8'b11111111;
memory[14578]=8'b11111111;
memory[14579]=8'b11111111;
memory[14580]=8'b11111111;
memory[14581]=8'b11111111;
memory[14582]=8'b11111111;
memory[14583]=8'b11111111;
memory[14584]=8'b00111111;
memory[14585]=8'b11111111;
memory[14586]=8'b11111111;
memory[14587]=8'b11111100;
memory[14588]=8'b01111111;
memory[14589]=8'b11111111;
memory[14590]=8'b11111111;
memory[14591]=8'b11111111;
memory[14592]=8'b11111111;
memory[14593]=8'b11111111;
memory[14594]=8'b11111111;
memory[14595]=8'b11111111;
memory[14596]=8'b11111111;
memory[14597]=8'b11111111;
memory[14598]=8'b11111111;
memory[14599]=8'b11111111;
memory[14600]=8'b11111111;
memory[14601]=8'b11111111;
memory[14602]=8'b11111111;
memory[14603]=8'b11111111;
memory[14604]=8'b11111111;
memory[14605]=8'b11111111;
memory[14606]=8'b11111111;
memory[14607]=8'b11111111;
memory[14608]=8'b11111111;
memory[14609]=8'b11111111;
memory[14610]=8'b11111111;
memory[14611]=8'b11111111;
memory[14612]=8'b11111111;
memory[14613]=8'b11111001;
memory[14614]=8'b11111111;
memory[14615]=8'b11111111;
memory[14616]=8'b11111111;
memory[14617]=8'b11111111;
memory[14618]=8'b11111111;
memory[14619]=8'b11111111;
memory[14620]=8'b11111111;
memory[14621]=8'b11111111;
memory[14622]=8'b11111111;
memory[14623]=8'b11111110;
memory[14624]=8'b01111111;
memory[14625]=8'b11100000;
memory[14626]=8'b00001111;
memory[14627]=8'b11111100;
memory[14628]=8'b11111111;
memory[14629]=8'b11111111;
memory[14630]=8'b11111111;
memory[14631]=8'b11111111;
memory[14632]=8'b11111111;
memory[14633]=8'b11111111;
memory[14634]=8'b11111111;
memory[14635]=8'b11111111;
memory[14636]=8'b11111111;
memory[14637]=8'b11111111;
memory[14638]=8'b11111111;
memory[14639]=8'b11111111;
memory[14640]=8'b11111111;
memory[14641]=8'b11111111;
memory[14642]=8'b11111111;
memory[14643]=8'b11111111;
memory[14644]=8'b11111111;
memory[14645]=8'b11111111;
memory[14646]=8'b11111111;
memory[14647]=8'b11111111;
memory[14648]=8'b11111111;
memory[14649]=8'b11111111;
memory[14650]=8'b11111111;
memory[14651]=8'b11111111;
memory[14652]=8'b11111111;
memory[14653]=8'b11111001;
memory[14654]=8'b11111111;
memory[14655]=8'b11111111;
memory[14656]=8'b11111111;
memory[14657]=8'b11111111;
memory[14658]=8'b11111111;
memory[14659]=8'b11111111;
memory[14660]=8'b11110001;
memory[14661]=8'b11111111;
memory[14662]=8'b11111111;
memory[14663]=8'b11110000;
memory[14664]=8'b11111111;
memory[14665]=8'b00001111;
memory[14666]=8'b11111111;
memory[14667]=8'b11111100;
memory[14668]=8'b11111111;
memory[14669]=8'b11111111;
memory[14670]=8'b11111111;
memory[14671]=8'b11111111;
memory[14672]=8'b11111111;
memory[14673]=8'b11111111;
memory[14674]=8'b11111111;
memory[14675]=8'b11111111;
memory[14676]=8'b11111111;
memory[14677]=8'b11111111;
memory[14678]=8'b11111111;
memory[14679]=8'b11111111;
memory[14680]=8'b11111111;
memory[14681]=8'b11111111;
memory[14682]=8'b11111111;
memory[14683]=8'b11111111;
memory[14684]=8'b11111111;
memory[14685]=8'b11111111;
memory[14686]=8'b11111111;
memory[14687]=8'b11111111;
memory[14688]=8'b11111111;
memory[14689]=8'b11111111;
memory[14690]=8'b11111111;
memory[14691]=8'b11111111;
memory[14692]=8'b11111111;
memory[14693]=8'b11011100;
memory[14694]=8'b11111111;
memory[14695]=8'b11111111;
memory[14696]=8'b11111111;
memory[14697]=8'b11111111;
memory[14698]=8'b11111111;
memory[14699]=8'b11111111;
memory[14700]=8'b11111111;
memory[14701]=8'b00000000;
memory[14702]=8'b00011100;
memory[14703]=8'b00000111;
memory[14704]=8'b11111000;
memory[14705]=8'b11111111;
memory[14706]=8'b11111111;
memory[14707]=8'b11111001;
memory[14708]=8'b11111111;
memory[14709]=8'b11111111;
memory[14710]=8'b11111111;
memory[14711]=8'b11111111;
memory[14712]=8'b11111111;
memory[14713]=8'b11111111;
memory[14714]=8'b11111111;
memory[14715]=8'b11111111;
memory[14716]=8'b11111111;
memory[14717]=8'b11111111;
memory[14718]=8'b11111111;
memory[14719]=8'b11111111;
memory[14720]=8'b11111111;
memory[14721]=8'b11111111;
memory[14722]=8'b11111111;
memory[14723]=8'b11111111;
memory[14724]=8'b11111111;
memory[14725]=8'b11111111;
memory[14726]=8'b11111111;
memory[14727]=8'b11111111;
memory[14728]=8'b11111111;
memory[14729]=8'b11111111;
memory[14730]=8'b11111111;
memory[14731]=8'b11111111;
memory[14732]=8'b11111111;
memory[14733]=8'b11001100;
memory[14734]=8'b11111111;
memory[14735]=8'b11111111;
memory[14736]=8'b11111111;
memory[14737]=8'b11111111;
memory[14738]=8'b11111111;
memory[14739]=8'b11111111;
memory[14740]=8'b11111111;
memory[14741]=8'b11111111;
memory[14742]=8'b10000011;
memory[14743]=8'b11111111;
memory[14744]=8'b10001111;
memory[14745]=8'b11111111;
memory[14746]=8'b11111111;
memory[14747]=8'b11111001;
memory[14748]=8'b11111111;
memory[14749]=8'b11111111;
memory[14750]=8'b11111111;
memory[14751]=8'b11111111;
memory[14752]=8'b11111111;
memory[14753]=8'b11111111;
memory[14754]=8'b11111111;
memory[14755]=8'b11111111;
memory[14756]=8'b11111111;
memory[14757]=8'b11111111;
memory[14758]=8'b11111111;
memory[14759]=8'b11111111;
memory[14760]=8'b11111111;
memory[14761]=8'b11111111;
memory[14762]=8'b11111111;
memory[14763]=8'b11111111;
memory[14764]=8'b11111111;
memory[14765]=8'b11111111;
memory[14766]=8'b11111111;
memory[14767]=8'b11111111;
memory[14768]=8'b11111111;
memory[14769]=8'b11111111;
memory[14770]=8'b11111111;
memory[14771]=8'b11111111;
memory[14772]=8'b11111111;
memory[14773]=8'b11001100;
memory[14774]=8'b11111111;
memory[14775]=8'b11111111;
memory[14776]=8'b11111111;
memory[14777]=8'b11111111;
memory[14778]=8'b11111111;
memory[14779]=8'b11111111;
memory[14780]=8'b11111111;
memory[14781]=8'b11111111;
memory[14782]=8'b11111111;
memory[14783]=8'b11111000;
memory[14784]=8'b11111111;
memory[14785]=8'b11111111;
memory[14786]=8'b11111111;
memory[14787]=8'b11111011;
memory[14788]=8'b11111111;
memory[14789]=8'b11111111;
memory[14790]=8'b11111111;
memory[14791]=8'b11111111;
memory[14792]=8'b11111111;
memory[14793]=8'b11111111;
memory[14794]=8'b11111111;
memory[14795]=8'b11111111;
memory[14796]=8'b11111111;
memory[14797]=8'b11111111;
memory[14798]=8'b11111111;
memory[14799]=8'b11111111;
memory[14800]=8'b11111111;
memory[14801]=8'b11111111;
memory[14802]=8'b11111111;
memory[14803]=8'b11111111;
memory[14804]=8'b11111111;
memory[14805]=8'b11111111;
memory[14806]=8'b11111111;
memory[14807]=8'b11111111;
memory[14808]=8'b11111111;
memory[14809]=8'b11111111;
memory[14810]=8'b11111111;
memory[14811]=8'b11111111;
memory[14812]=8'b11111111;
memory[14813]=8'b11101100;
memory[14814]=8'b01111111;
memory[14815]=8'b11111111;
memory[14816]=8'b11111111;
memory[14817]=8'b11111111;
memory[14818]=8'b11111111;
memory[14819]=8'b11111111;
memory[14820]=8'b11111111;
memory[14821]=8'b11111111;
memory[14822]=8'b11111111;
memory[14823]=8'b11111111;
memory[14824]=8'b11111111;
memory[14825]=8'b11111111;
memory[14826]=8'b11111111;
memory[14827]=8'b11111011;
memory[14828]=8'b11111111;
memory[14829]=8'b11111001;
memory[14830]=8'b11111111;
memory[14831]=8'b11111111;
memory[14832]=8'b11111111;
memory[14833]=8'b11111111;
memory[14834]=8'b11111111;
memory[14835]=8'b11111111;
memory[14836]=8'b11111111;
memory[14837]=8'b11111111;
memory[14838]=8'b11111111;
memory[14839]=8'b11111111;
memory[14840]=8'b11111111;
memory[14841]=8'b11111111;
memory[14842]=8'b11111111;
memory[14843]=8'b11111111;
memory[14844]=8'b11111111;
memory[14845]=8'b11111111;
memory[14846]=8'b11111111;
memory[14847]=8'b11111111;
memory[14848]=8'b11111111;
memory[14849]=8'b11111111;
memory[14850]=8'b11111111;
memory[14851]=8'b11111111;
memory[14852]=8'b11111111;
memory[14853]=8'b11001100;
memory[14854]=8'b01111111;
memory[14855]=8'b11111111;
memory[14856]=8'b11111111;
memory[14857]=8'b00000000;
memory[14858]=8'b00000111;
memory[14859]=8'b11111111;
memory[14860]=8'b11111111;
memory[14861]=8'b11111111;
memory[14862]=8'b11111111;
memory[14863]=8'b11111111;
memory[14864]=8'b11111111;
memory[14865]=8'b11111111;
memory[14866]=8'b11111111;
memory[14867]=8'b11110011;
memory[14868]=8'b11111111;
memory[14869]=8'b11000000;
memory[14870]=8'b00011111;
memory[14871]=8'b11111111;
memory[14872]=8'b11111111;
memory[14873]=8'b11111111;
memory[14874]=8'b11111111;
memory[14875]=8'b11111111;
memory[14876]=8'b11111111;
memory[14877]=8'b11111111;
memory[14878]=8'b11111111;
memory[14879]=8'b11111111;
memory[14880]=8'b11111111;
memory[14881]=8'b11111111;
memory[14882]=8'b11111111;
memory[14883]=8'b11111111;
memory[14884]=8'b11111111;
memory[14885]=8'b11111111;
memory[14886]=8'b11111111;
memory[14887]=8'b11111111;
memory[14888]=8'b11111111;
memory[14889]=8'b11111111;
memory[14890]=8'b11111111;
memory[14891]=8'b11111111;
memory[14892]=8'b11111111;
memory[14893]=8'b11000110;
memory[14894]=8'b01111111;
memory[14895]=8'b11111111;
memory[14896]=8'b11111111;
memory[14897]=8'b11111110;
memory[14898]=8'b00000000;
memory[14899]=8'b00000111;
memory[14900]=8'b11111111;
memory[14901]=8'b11111111;
memory[14902]=8'b11111111;
memory[14903]=8'b11111111;
memory[14904]=8'b11111111;
memory[14905]=8'b11111111;
memory[14906]=8'b11111111;
memory[14907]=8'b11110001;
memory[14908]=8'b11111111;
memory[14909]=8'b11111111;
memory[14910]=8'b00000011;
memory[14911]=8'b11111111;
memory[14912]=8'b11111111;
memory[14913]=8'b11111111;
memory[14914]=8'b11111111;
memory[14915]=8'b11111111;
memory[14916]=8'b11111111;
memory[14917]=8'b11111111;
memory[14918]=8'b11111111;
memory[14919]=8'b11111111;
memory[14920]=8'b11111111;
memory[14921]=8'b11111111;
memory[14922]=8'b11111111;
memory[14923]=8'b11111111;
memory[14924]=8'b11111111;
memory[14925]=8'b11111111;
memory[14926]=8'b11111111;
memory[14927]=8'b11111000;
memory[14928]=8'b00000000;
memory[14929]=8'b11111111;
memory[14930]=8'b11111111;
memory[14931]=8'b11111111;
memory[14932]=8'b11111111;
memory[14933]=8'b11100010;
memory[14934]=8'b00111111;
memory[14935]=8'b11111111;
memory[14936]=8'b11111111;
memory[14937]=8'b11111111;
memory[14938]=8'b11111000;
memory[14939]=8'b00000000;
memory[14940]=8'b01111111;
memory[14941]=8'b11111111;
memory[14942]=8'b11111111;
memory[14943]=8'b11111111;
memory[14944]=8'b00011111;
memory[14945]=8'b11111111;
memory[14946]=8'b11111111;
memory[14947]=8'b11110001;
memory[14948]=8'b11111111;
memory[14949]=8'b11111111;
memory[14950]=8'b11110000;
memory[14951]=8'b00000000;
memory[14952]=8'b11111111;
memory[14953]=8'b11111111;
memory[14954]=8'b11111111;
memory[14955]=8'b11111111;
memory[14956]=8'b11111111;
memory[14957]=8'b11111111;
memory[14958]=8'b11111111;
memory[14959]=8'b11111111;
memory[14960]=8'b11111111;
memory[14961]=8'b11111111;
memory[14962]=8'b11111111;
memory[14963]=8'b11111111;
memory[14964]=8'b11111111;
memory[14965]=8'b11111111;
memory[14966]=8'b11111111;
memory[14967]=8'b11111111;
memory[14968]=8'b11111100;
memory[14969]=8'b00001111;
memory[14970]=8'b11111111;
memory[14971]=8'b11111111;
memory[14972]=8'b11111111;
memory[14973]=8'b11000011;
memory[14974]=8'b00111111;
memory[14975]=8'b11111111;
memory[14976]=8'b11111111;
memory[14977]=8'b11111111;
memory[14978]=8'b11111111;
memory[14979]=8'b10000000;
memory[14980]=8'b00000111;
memory[14981]=8'b11111111;
memory[14982]=8'b11111111;
memory[14983]=8'b11100000;
memory[14984]=8'b11111111;
memory[14985]=8'b11111111;
memory[14986]=8'b11111111;
memory[14987]=8'b11100101;
memory[14988]=8'b11111111;
memory[14989]=8'b11111111;
memory[14990]=8'b11111111;
memory[14991]=8'b11111111;
memory[14992]=8'b11111111;
memory[14993]=8'b11111111;
memory[14994]=8'b11111111;
memory[14995]=8'b11111111;
memory[14996]=8'b11111111;
memory[14997]=8'b11111111;
memory[14998]=8'b11111111;
memory[14999]=8'b11111111;
memory[15000]=8'b11111111;
memory[15001]=8'b11111111;
memory[15002]=8'b11111111;
memory[15003]=8'b11111111;
memory[15004]=8'b11111111;
memory[15005]=8'b11111111;
memory[15006]=8'b11111111;
memory[15007]=8'b11111111;
memory[15008]=8'b11111111;
memory[15009]=8'b11000001;
memory[15010]=8'b11111111;
memory[15011]=8'b11111111;
memory[15012]=8'b11111111;
memory[15013]=8'b11000011;
memory[15014]=8'b00111111;
memory[15015]=8'b11111111;
memory[15016]=8'b11111111;
memory[15017]=8'b11111111;
memory[15018]=8'b11111111;
memory[15019]=8'b11111000;
memory[15020]=8'b00000000;
memory[15021]=8'b00111111;
memory[15022]=8'b11000000;
memory[15023]=8'b00000111;
memory[15024]=8'b11111111;
memory[15025]=8'b11111111;
memory[15026]=8'b11111111;
memory[15027]=8'b11100001;
memory[15028]=8'b11111111;
memory[15029]=8'b11111111;
memory[15030]=8'b11111111;
memory[15031]=8'b11111111;
memory[15032]=8'b11111111;
memory[15033]=8'b11111111;
memory[15034]=8'b11111111;
memory[15035]=8'b11111111;
memory[15036]=8'b11111111;
memory[15037]=8'b11111111;
memory[15038]=8'b11111111;
memory[15039]=8'b11111111;
memory[15040]=8'b11111111;
memory[15041]=8'b11111111;
memory[15042]=8'b11111111;
memory[15043]=8'b11111111;
memory[15044]=8'b11111111;
memory[15045]=8'b11111111;
memory[15046]=8'b11111111;
memory[15047]=8'b11111111;
memory[15048]=8'b11111111;
memory[15049]=8'b11110000;
memory[15050]=8'b00111111;
memory[15051]=8'b10111111;
memory[15052]=8'b11111111;
memory[15053]=8'b11000011;
memory[15054]=8'b00011111;
memory[15055]=8'b11111111;
memory[15056]=8'b11111111;
memory[15057]=8'b11111111;
memory[15058]=8'b11111111;
memory[15059]=8'b11111111;
memory[15060]=8'b10000000;
memory[15061]=8'b00000000;
memory[15062]=8'b00000000;
memory[15063]=8'b01111111;
memory[15064]=8'b11111111;
memory[15065]=8'b11111111;
memory[15066]=8'b11111111;
memory[15067]=8'b11100001;
memory[15068]=8'b11111111;
memory[15069]=8'b11111111;
memory[15070]=8'b11111111;
memory[15071]=8'b11111111;
memory[15072]=8'b11111111;
memory[15073]=8'b11111111;
memory[15074]=8'b11111111;
memory[15075]=8'b11111111;
memory[15076]=8'b11111111;
memory[15077]=8'b11111111;
memory[15078]=8'b11111111;
memory[15079]=8'b11111111;
memory[15080]=8'b11111111;
memory[15081]=8'b11111111;
memory[15082]=8'b11111111;
memory[15083]=8'b11111111;
memory[15084]=8'b11111111;
memory[15085]=8'b11111111;
memory[15086]=8'b11111111;
memory[15087]=8'b11111111;
memory[15088]=8'b11111111;
memory[15089]=8'b11111111;
memory[15090]=8'b10000111;
memory[15091]=8'b11111111;
memory[15092]=8'b11111111;
memory[15093]=8'b11000011;
memory[15094]=8'b00011111;
memory[15095]=8'b11111111;
memory[15096]=8'b11111111;
memory[15097]=8'b11111111;
memory[15098]=8'b11111111;
memory[15099]=8'b11111111;
memory[15100]=8'b11111111;
memory[15101]=8'b10000001;
memory[15102]=8'b11111111;
memory[15103]=8'b11111111;
memory[15104]=8'b11111111;
memory[15105]=8'b11111111;
memory[15106]=8'b11111111;
memory[15107]=8'b11100001;
memory[15108]=8'b11111111;
memory[15109]=8'b11111111;
memory[15110]=8'b11111111;
memory[15111]=8'b11111111;
memory[15112]=8'b11111111;
memory[15113]=8'b11111111;
memory[15114]=8'b11111111;
memory[15115]=8'b11111111;
memory[15116]=8'b11111111;
memory[15117]=8'b11111111;
memory[15118]=8'b11111111;
memory[15119]=8'b11111111;
memory[15120]=8'b11111111;
memory[15121]=8'b11111111;
memory[15122]=8'b11111111;
memory[15123]=8'b11111111;
memory[15124]=8'b11111111;
memory[15125]=8'b11111111;
memory[15126]=8'b11111111;
memory[15127]=8'b11111111;
memory[15128]=8'b11111111;
memory[15129]=8'b11111111;
memory[15130]=8'b11111111;
memory[15131]=8'b11111111;
memory[15132]=8'b11111111;
memory[15133]=8'b11000011;
memory[15134]=8'b00011111;
memory[15135]=8'b11111111;
memory[15136]=8'b11111111;
memory[15137]=8'b11111111;
memory[15138]=8'b11111111;
memory[15139]=8'b11111111;
memory[15140]=8'b11111111;
memory[15141]=8'b11111111;
memory[15142]=8'b11111111;
memory[15143]=8'b11111111;
memory[15144]=8'b11111111;
memory[15145]=8'b11111111;
memory[15146]=8'b11111111;
memory[15147]=8'b11000001;
memory[15148]=8'b11111111;
memory[15149]=8'b11111111;
memory[15150]=8'b11111111;
memory[15151]=8'b11111111;
memory[15152]=8'b11111111;
memory[15153]=8'b11111111;
memory[15154]=8'b11111111;
memory[15155]=8'b11111111;
memory[15156]=8'b11111111;
memory[15157]=8'b11111111;
memory[15158]=8'b11111111;
memory[15159]=8'b11111111;
memory[15160]=8'b11111111;
memory[15161]=8'b11111111;
memory[15162]=8'b11111111;
memory[15163]=8'b11111111;
memory[15164]=8'b11111111;
memory[15165]=8'b11111111;
memory[15166]=8'b11111111;
memory[15167]=8'b11111111;
memory[15168]=8'b11111111;
memory[15169]=8'b11111111;
memory[15170]=8'b11111111;
memory[15171]=8'b11111111;
memory[15172]=8'b11111111;
memory[15173]=8'b11000111;
memory[15174]=8'b00011111;
memory[15175]=8'b11111111;
memory[15176]=8'b11111111;
memory[15177]=8'b11111111;
memory[15178]=8'b11111111;
memory[15179]=8'b11111111;
memory[15180]=8'b11111111;
memory[15181]=8'b11111111;
memory[15182]=8'b11111111;
memory[15183]=8'b11111111;
memory[15184]=8'b11111111;
memory[15185]=8'b11111111;
memory[15186]=8'b11111111;
memory[15187]=8'b11001001;
memory[15188]=8'b11111111;
memory[15189]=8'b11111111;
memory[15190]=8'b11111111;
memory[15191]=8'b11111111;
memory[15192]=8'b11111111;
memory[15193]=8'b11111111;
memory[15194]=8'b11111111;
memory[15195]=8'b11111111;
memory[15196]=8'b11111111;
memory[15197]=8'b11111111;
memory[15198]=8'b11111111;
memory[15199]=8'b11111111;
memory[15200]=8'b11111111;
memory[15201]=8'b11111111;
memory[15202]=8'b11111111;
memory[15203]=8'b11111111;
memory[15204]=8'b11111111;
memory[15205]=8'b11111111;
memory[15206]=8'b11111111;
memory[15207]=8'b11111111;
memory[15208]=8'b11111111;
memory[15209]=8'b11111111;
memory[15210]=8'b11111111;
memory[15211]=8'b11111111;
memory[15212]=8'b11111111;
memory[15213]=8'b11000011;
memory[15214]=8'b00001111;
memory[15215]=8'b11111111;
memory[15216]=8'b11111111;
memory[15217]=8'b11111111;
memory[15218]=8'b11111111;
memory[15219]=8'b11111111;
memory[15220]=8'b11111111;
memory[15221]=8'b11111111;
memory[15222]=8'b11111111;
memory[15223]=8'b11111111;
memory[15224]=8'b11111111;
memory[15225]=8'b11111111;
memory[15226]=8'b11111111;
memory[15227]=8'b11001001;
memory[15228]=8'b11111111;
memory[15229]=8'b11111111;
memory[15230]=8'b11111111;
memory[15231]=8'b11111111;
memory[15232]=8'b11111111;
memory[15233]=8'b11111111;
memory[15234]=8'b11111111;
memory[15235]=8'b11111111;
memory[15236]=8'b11111111;
memory[15237]=8'b11111111;
memory[15238]=8'b11111111;
memory[15239]=8'b11111111;
memory[15240]=8'b11111111;
memory[15241]=8'b11111111;
memory[15242]=8'b11111111;
memory[15243]=8'b11111111;
memory[15244]=8'b11111111;
memory[15245]=8'b11111111;
memory[15246]=8'b11111111;
memory[15247]=8'b11111111;
memory[15248]=8'b11111111;
memory[15249]=8'b11111111;
memory[15250]=8'b11111111;
memory[15251]=8'b11111111;
memory[15252]=8'b11111111;
memory[15253]=8'b11000011;
memory[15254]=8'b00000111;
memory[15255]=8'b11111111;
memory[15256]=8'b11111111;
memory[15257]=8'b11111111;
memory[15258]=8'b11111111;
memory[15259]=8'b11111111;
memory[15260]=8'b11111111;
memory[15261]=8'b11111111;
memory[15262]=8'b11111111;
memory[15263]=8'b11111111;
memory[15264]=8'b11111111;
memory[15265]=8'b11111111;
memory[15266]=8'b11111111;
memory[15267]=8'b10011001;
memory[15268]=8'b11111111;
memory[15269]=8'b11111111;
memory[15270]=8'b11111111;
memory[15271]=8'b11111111;
memory[15272]=8'b11111111;
memory[15273]=8'b11111111;
memory[15274]=8'b11111111;
memory[15275]=8'b11111111;
memory[15276]=8'b11111111;
memory[15277]=8'b11111111;
memory[15278]=8'b11111111;
memory[15279]=8'b11111111;
memory[15280]=8'b11111111;
memory[15281]=8'b11111111;
memory[15282]=8'b11111111;
memory[15283]=8'b11111111;
memory[15284]=8'b11111111;
memory[15285]=8'b11111111;
memory[15286]=8'b11111111;
memory[15287]=8'b11111111;
memory[15288]=8'b11111111;
memory[15289]=8'b11111111;
memory[15290]=8'b11111111;
memory[15291]=8'b11111111;
memory[15292]=8'b11111111;
memory[15293]=8'b10000001;
memory[15294]=8'b00000111;
memory[15295]=8'b11111111;
memory[15296]=8'b11111111;
memory[15297]=8'b11111111;
memory[15298]=8'b11111111;
memory[15299]=8'b11111111;
memory[15300]=8'b11111111;
memory[15301]=8'b11111111;
memory[15302]=8'b11111111;
memory[15303]=8'b11111111;
memory[15304]=8'b11111111;
memory[15305]=8'b11111111;
memory[15306]=8'b11111111;
memory[15307]=8'b10011001;
memory[15308]=8'b11111111;
memory[15309]=8'b11111111;
memory[15310]=8'b11111111;
memory[15311]=8'b11111111;
memory[15312]=8'b11111111;
memory[15313]=8'b11111111;
memory[15314]=8'b11111111;
memory[15315]=8'b11111111;
memory[15316]=8'b11111111;
memory[15317]=8'b11111111;
memory[15318]=8'b11111111;
memory[15319]=8'b11111111;
memory[15320]=8'b11111111;
memory[15321]=8'b11111111;
memory[15322]=8'b11111111;
memory[15323]=8'b11111111;
memory[15324]=8'b11111111;
memory[15325]=8'b11111111;
memory[15326]=8'b11111111;
memory[15327]=8'b11111111;
memory[15328]=8'b11111111;
memory[15329]=8'b11111111;
memory[15330]=8'b11111111;
memory[15331]=8'b11111111;
memory[15332]=8'b11111111;
memory[15333]=8'b10000001;
memory[15334]=8'b10000001;
memory[15335]=8'b11111111;
memory[15336]=8'b11111111;
memory[15337]=8'b11111111;
memory[15338]=8'b11111111;
memory[15339]=8'b11111111;
memory[15340]=8'b11111111;
memory[15341]=8'b11111111;
memory[15342]=8'b11111111;
memory[15343]=8'b11111111;
memory[15344]=8'b11111111;
memory[15345]=8'b11111111;
memory[15346]=8'b11111111;
memory[15347]=8'b10011001;
memory[15348]=8'b11111111;
memory[15349]=8'b11111111;
memory[15350]=8'b11111111;
memory[15351]=8'b11111111;
memory[15352]=8'b11111111;
memory[15353]=8'b11111111;
memory[15354]=8'b11111111;
memory[15355]=8'b11111111;
memory[15356]=8'b11111111;
memory[15357]=8'b11111111;
memory[15358]=8'b11111111;
memory[15359]=8'b11111111;
memory[15360]=8'b11111111;
memory[15361]=8'b11111111;
memory[15362]=8'b11111111;
memory[15363]=8'b11111111;
memory[15364]=8'b11111111;
memory[15365]=8'b11111111;
memory[15366]=8'b11111111;
memory[15367]=8'b11111111;
memory[15368]=8'b11111111;
memory[15369]=8'b11111111;
memory[15370]=8'b11111111;
memory[15371]=8'b11111111;
memory[15372]=8'b11111111;
memory[15373]=8'b00000001;
memory[15374]=8'b10000000;
memory[15375]=8'b00111111;
memory[15376]=8'b11111111;
memory[15377]=8'b11111111;
memory[15378]=8'b11111111;
memory[15379]=8'b11111111;
memory[15380]=8'b11111111;
memory[15381]=8'b11111111;
memory[15382]=8'b11111111;
memory[15383]=8'b11111111;
memory[15384]=8'b11111111;
memory[15385]=8'b11111111;
memory[15386]=8'b11111111;
memory[15387]=8'b00011000;
memory[15388]=8'b11111111;
memory[15389]=8'b11111111;
memory[15390]=8'b11111111;
memory[15391]=8'b11111111;
memory[15392]=8'b11111111;
memory[15393]=8'b11111111;
memory[15394]=8'b11111111;
memory[15395]=8'b11111111;
memory[15396]=8'b11111111;
memory[15397]=8'b11111111;
memory[15398]=8'b11111111;
memory[15399]=8'b11111111;
memory[15400]=8'b11111111;
memory[15401]=8'b11111111;
memory[15402]=8'b11111111;
memory[15403]=8'b11111111;
memory[15404]=8'b11111111;
memory[15405]=8'b11111111;
memory[15406]=8'b11111111;
memory[15407]=8'b11111111;
memory[15408]=8'b11111111;
memory[15409]=8'b11111111;
memory[15410]=8'b11111111;
memory[15411]=8'b11111111;
memory[15412]=8'b11111110;
memory[15413]=8'b00000000;
memory[15414]=8'b11000000;
memory[15415]=8'b00000111;
memory[15416]=8'b11111111;
memory[15417]=8'b11111111;
memory[15418]=8'b11111111;
memory[15419]=8'b11111111;
memory[15420]=8'b11111111;
memory[15421]=8'b11111111;
memory[15422]=8'b11111111;
memory[15423]=8'b11111111;
memory[15424]=8'b11111111;
memory[15425]=8'b11111111;
memory[15426]=8'b11111110;
memory[15427]=8'b00000000;
memory[15428]=8'b11111111;
memory[15429]=8'b11111111;
memory[15430]=8'b11111111;
memory[15431]=8'b11111111;
memory[15432]=8'b11111111;
memory[15433]=8'b11111111;
memory[15434]=8'b11111111;
memory[15435]=8'b11111111;
memory[15436]=8'b11111111;
memory[15437]=8'b11111111;
memory[15438]=8'b11111111;
memory[15439]=8'b11111111;
memory[15440]=8'b11111111;
memory[15441]=8'b11111111;
memory[15442]=8'b11111111;
memory[15443]=8'b11111111;
memory[15444]=8'b11111111;
memory[15445]=8'b11111111;
memory[15446]=8'b11111111;
memory[15447]=8'b11111111;
memory[15448]=8'b11111111;
memory[15449]=8'b11111111;
memory[15450]=8'b11111111;
memory[15451]=8'b11111111;
memory[15452]=8'b11111100;
memory[15453]=8'b00000000;
memory[15454]=8'b11000000;
memory[15455]=8'b00000000;
memory[15456]=8'b11111111;
memory[15457]=8'b11111111;
memory[15458]=8'b11111111;
memory[15459]=8'b11111111;
memory[15460]=8'b11111111;
memory[15461]=8'b11111111;
memory[15462]=8'b11111111;
memory[15463]=8'b11111111;
memory[15464]=8'b11111111;
memory[15465]=8'b11111111;
memory[15466]=8'b11111100;
memory[15467]=8'b00000000;
memory[15468]=8'b01111111;
memory[15469]=8'b11111111;
memory[15470]=8'b11111111;
memory[15471]=8'b11111111;
memory[15472]=8'b11111111;
memory[15473]=8'b11111111;
memory[15474]=8'b11111111;
memory[15475]=8'b11111111;
memory[15476]=8'b11111111;
memory[15477]=8'b11111111;
memory[15478]=8'b11111111;
memory[15479]=8'b11111111;
memory[15480]=8'b11111111;
memory[15481]=8'b11111111;
memory[15482]=8'b11111111;
memory[15483]=8'b11111111;
memory[15484]=8'b11111111;
memory[15485]=8'b11111111;
memory[15486]=8'b11111111;
memory[15487]=8'b11111111;
memory[15488]=8'b11111111;
memory[15489]=8'b11111111;
memory[15490]=8'b11111111;
memory[15491]=8'b11111111;
memory[15492]=8'b11111111;
memory[15493]=8'b11111111;
memory[15494]=8'b11100000;
memory[15495]=8'b00000000;
memory[15496]=8'b00001111;
memory[15497]=8'b11111111;
memory[15498]=8'b11111111;
memory[15499]=8'b11111111;
memory[15500]=8'b11111111;
memory[15501]=8'b11111111;
memory[15502]=8'b11111111;
memory[15503]=8'b11111111;
memory[15504]=8'b11111111;
memory[15505]=8'b11111111;
memory[15506]=8'b11100000;
memory[15507]=8'b00000000;
memory[15508]=8'b00111111;
memory[15509]=8'b11111111;
memory[15510]=8'b11111111;
memory[15511]=8'b11111111;
memory[15512]=8'b11111111;
memory[15513]=8'b11111111;
memory[15514]=8'b11111111;
memory[15515]=8'b11111111;
memory[15516]=8'b11111111;
memory[15517]=8'b11111111;
memory[15518]=8'b11111111;
memory[15519]=8'b11111111;
memory[15520]=8'b11111111;
memory[15521]=8'b11111111;
memory[15522]=8'b11111111;
memory[15523]=8'b11111111;
memory[15524]=8'b11111111;
memory[15525]=8'b11111111;
memory[15526]=8'b11111111;
memory[15527]=8'b11111111;
memory[15528]=8'b11111111;
memory[15529]=8'b11111111;
memory[15530]=8'b11111111;
memory[15531]=8'b11111111;
memory[15532]=8'b11111111;
memory[15533]=8'b11111111;
memory[15534]=8'b11100111;
memory[15535]=8'b10000000;
memory[15536]=8'b00000001;
memory[15537]=8'b11111111;
memory[15538]=8'b11111111;
memory[15539]=8'b11111111;
memory[15540]=8'b11111111;
memory[15541]=8'b11111111;
memory[15542]=8'b11111111;
memory[15543]=8'b11111111;
memory[15544]=8'b11111111;
memory[15545]=8'b11111110;
memory[15546]=8'b00000000;
memory[15547]=8'b00110000;
memory[15548]=8'b00111111;
memory[15549]=8'b11111111;
memory[15550]=8'b11111111;
memory[15551]=8'b11111111;
memory[15552]=8'b11111111;
memory[15553]=8'b11111111;
memory[15554]=8'b11111111;
memory[15555]=8'b11111111;
memory[15556]=8'b11111111;
memory[15557]=8'b11111111;
memory[15558]=8'b11111111;
memory[15559]=8'b11111111;
memory[15560]=8'b11111111;
memory[15561]=8'b11111111;
memory[15562]=8'b11111111;
memory[15563]=8'b11111111;
memory[15564]=8'b11111111;
memory[15565]=8'b11111111;
memory[15566]=8'b11111111;
memory[15567]=8'b11111111;
memory[15568]=8'b11111111;
memory[15569]=8'b11111111;
memory[15570]=8'b11111111;
memory[15571]=8'b11111111;
memory[15572]=8'b11111111;
memory[15573]=8'b11111111;
memory[15574]=8'b11111111;
memory[15575]=8'b11111111;
memory[15576]=8'b11111111;
memory[15577]=8'b11111111;
memory[15578]=8'b11111111;
memory[15579]=8'b11111111;
memory[15580]=8'b11111111;
memory[15581]=8'b11111111;
memory[15582]=8'b11111111;
memory[15583]=8'b11111111;
memory[15584]=8'b11111111;
memory[15585]=8'b11100000;
memory[15586]=8'b00000000;
memory[15587]=8'b01111111;
memory[15588]=8'b11111111;
memory[15589]=8'b11111111;
memory[15590]=8'b11111111;
memory[15591]=8'b11111111;
memory[15592]=8'b11111111;
memory[15593]=8'b11111111;
memory[15594]=8'b11111111;
memory[15595]=8'b11111111;
memory[15596]=8'b11111111;
memory[15597]=8'b11111111;
memory[15598]=8'b11111111;
memory[15599]=8'b11111111;
memory[15600]=8'b11111111;
memory[15601]=8'b11111111;
memory[15602]=8'b11111111;
memory[15603]=8'b11111111;
memory[15604]=8'b11111111;
memory[15605]=8'b11111111;
memory[15606]=8'b11111111;
memory[15607]=8'b11111111;
memory[15608]=8'b11111111;
memory[15609]=8'b11111111;
memory[15610]=8'b11111111;
memory[15611]=8'b11111111;
memory[15612]=8'b11111111;
memory[15613]=8'b11111111;
memory[15614]=8'b11111111;
memory[15615]=8'b11111111;
memory[15616]=8'b11111111;
memory[15617]=8'b11111111;
memory[15618]=8'b11111111;
memory[15619]=8'b11111111;
memory[15620]=8'b11111111;
memory[15621]=8'b11111111;
memory[15622]=8'b11111111;
memory[15623]=8'b11111111;
memory[15624]=8'b11111111;
memory[15625]=8'b11111111;
memory[15626]=8'b11111111;
memory[15627]=8'b11111111;
memory[15628]=8'b11111111;
memory[15629]=8'b11111111;
memory[15630]=8'b11111111;
memory[15631]=8'b11111111;
memory[15632]=8'b11111111;
memory[15633]=8'b11111111;
memory[15634]=8'b11111111;
memory[15635]=8'b11111111;
memory[15636]=8'b11111111;
memory[15637]=8'b11111111;
memory[15638]=8'b11111111;
memory[15639]=8'b11111111;
memory[15640]=8'b11111111;
memory[15641]=8'b11111111;
memory[15642]=8'b11111111;
memory[15643]=8'b11111111;
memory[15644]=8'b11111111;
memory[15645]=8'b11111111;
memory[15646]=8'b11111111;
memory[15647]=8'b11111111;
memory[15648]=8'b11111111;
memory[15649]=8'b11111111;
memory[15650]=8'b11111111;
memory[15651]=8'b11111111;
memory[15652]=8'b11111111;
memory[15653]=8'b11111111;
memory[15654]=8'b11111111;
memory[15655]=8'b11111111;
memory[15656]=8'b11111111;
memory[15657]=8'b11111111;
memory[15658]=8'b11111111;
memory[15659]=8'b11111111;
memory[15660]=8'b11111111;
memory[15661]=8'b11111111;
memory[15662]=8'b11111111;
memory[15663]=8'b11111111;
memory[15664]=8'b11111111;
memory[15665]=8'b11111111;
memory[15666]=8'b11111111;
memory[15667]=8'b11111111;
memory[15668]=8'b11111111;
memory[15669]=8'b11111111;
memory[15670]=8'b11111111;
memory[15671]=8'b11111111;
memory[15672]=8'b11111111;
memory[15673]=8'b11111111;
memory[15674]=8'b11111111;
memory[15675]=8'b11111111;
memory[15676]=8'b11111111;
memory[15677]=8'b11111111;
memory[15678]=8'b11111111;
memory[15679]=8'b11111111;
memory[15680]=8'b11111111;
memory[15681]=8'b11111111;
memory[15682]=8'b11111111;
memory[15683]=8'b11111111;
memory[15684]=8'b11111111;
memory[15685]=8'b11111111;
memory[15686]=8'b11111111;
memory[15687]=8'b11111111;
memory[15688]=8'b11111111;
memory[15689]=8'b11111111;
memory[15690]=8'b11111111;
memory[15691]=8'b11111111;
memory[15692]=8'b11111111;
memory[15693]=8'b11111111;
memory[15694]=8'b11111111;
memory[15695]=8'b11111111;
memory[15696]=8'b11111111;
memory[15697]=8'b11111111;
memory[15698]=8'b11111111;
memory[15699]=8'b11111111;
memory[15700]=8'b11111111;
memory[15701]=8'b11111111;
memory[15702]=8'b11111111;
memory[15703]=8'b11111111;
memory[15704]=8'b11111111;
memory[15705]=8'b11111111;
memory[15706]=8'b11111111;
memory[15707]=8'b11111111;
memory[15708]=8'b11111111;
memory[15709]=8'b11111111;
memory[15710]=8'b11111111;
memory[15711]=8'b11111111;
memory[15712]=8'b11111111;
memory[15713]=8'b11111111;
memory[15714]=8'b11111111;
memory[15715]=8'b11111111;
memory[15716]=8'b11111111;
memory[15717]=8'b11111111;
memory[15718]=8'b11111111;
memory[15719]=8'b11111111;
memory[15720]=8'b11111111;
memory[15721]=8'b11111111;
memory[15722]=8'b11111111;
memory[15723]=8'b11111111;
memory[15724]=8'b11111111;
memory[15725]=8'b11111111;
memory[15726]=8'b11111111;
memory[15727]=8'b11111111;
memory[15728]=8'b11111111;
memory[15729]=8'b11111111;
memory[15730]=8'b11111111;
memory[15731]=8'b11111111;
memory[15732]=8'b11111111;
memory[15733]=8'b11111111;
memory[15734]=8'b11111111;
memory[15735]=8'b11111111;
memory[15736]=8'b11111111;
memory[15737]=8'b11111111;
memory[15738]=8'b11111111;
memory[15739]=8'b11111111;
memory[15740]=8'b11111111;
memory[15741]=8'b11111111;
memory[15742]=8'b11111111;
memory[15743]=8'b11111111;
memory[15744]=8'b11111111;
memory[15745]=8'b11111111;
memory[15746]=8'b11111111;
memory[15747]=8'b11111111;
memory[15748]=8'b11111111;
memory[15749]=8'b11111111;
memory[15750]=8'b11111111;
memory[15751]=8'b11111111;
memory[15752]=8'b11111111;
memory[15753]=8'b11111111;
memory[15754]=8'b11111111;
memory[15755]=8'b11111111;
memory[15756]=8'b11111111;
memory[15757]=8'b11111111;
memory[15758]=8'b11111111;
memory[15759]=8'b11111111;
memory[15760]=8'b11111111;
memory[15761]=8'b11111111;
memory[15762]=8'b11111111;
memory[15763]=8'b11111111;
memory[15764]=8'b11111111;
memory[15765]=8'b11111111;
memory[15766]=8'b11111111;
memory[15767]=8'b11111111;
memory[15768]=8'b11111111;
memory[15769]=8'b11111111;
memory[15770]=8'b11111111;
memory[15771]=8'b11111111;
memory[15772]=8'b11111111;
memory[15773]=8'b11111111;
memory[15774]=8'b11111111;
memory[15775]=8'b11111111;
memory[15776]=8'b11111111;
memory[15777]=8'b11111111;
memory[15778]=8'b11111111;
memory[15779]=8'b11111111;
memory[15780]=8'b11111111;
memory[15781]=8'b11111111;
memory[15782]=8'b11111111;
memory[15783]=8'b11111111;
memory[15784]=8'b11111111;
memory[15785]=8'b11111111;
memory[15786]=8'b11111111;
memory[15787]=8'b11111111;
memory[15788]=8'b11111111;
memory[15789]=8'b11111111;
memory[15790]=8'b11111111;
memory[15791]=8'b11111111;
memory[15792]=8'b11111111;
memory[15793]=8'b11111111;
memory[15794]=8'b11111111;
memory[15795]=8'b11111111;
memory[15796]=8'b11111111;
memory[15797]=8'b11111111;
memory[15798]=8'b11111111;
memory[15799]=8'b11111111;
memory[15800]=8'b11111111;
memory[15801]=8'b11111111;
memory[15802]=8'b11111111;
memory[15803]=8'b11111111;
memory[15804]=8'b11111111;
memory[15805]=8'b11111111;
memory[15806]=8'b11111111;
memory[15807]=8'b11111111;
memory[15808]=8'b11111111;
memory[15809]=8'b11111111;
memory[15810]=8'b11111111;
memory[15811]=8'b11111111;
memory[15812]=8'b11111111;
memory[15813]=8'b11111111;
memory[15814]=8'b11111111;
memory[15815]=8'b11111111;
memory[15816]=8'b11111111;
memory[15817]=8'b11111111;
memory[15818]=8'b11111111;
memory[15819]=8'b11111111;
memory[15820]=8'b11111111;
memory[15821]=8'b11111111;
memory[15822]=8'b11111111;
memory[15823]=8'b11111111;
memory[15824]=8'b11111111;
memory[15825]=8'b11111111;
memory[15826]=8'b11111111;
memory[15827]=8'b11111111;
memory[15828]=8'b11111111;
memory[15829]=8'b11111111;
memory[15830]=8'b11111111;
memory[15831]=8'b11111111;
memory[15832]=8'b11111111;
memory[15833]=8'b11111111;
memory[15834]=8'b11111111;
memory[15835]=8'b11111111;
memory[15836]=8'b11111111;
memory[15837]=8'b11111111;
memory[15838]=8'b11111111;
memory[15839]=8'b11111111;
memory[15840]=8'b11111111;
memory[15841]=8'b11111111;
memory[15842]=8'b11111111;
memory[15843]=8'b11111111;
memory[15844]=8'b11111111;
memory[15845]=8'b11111111;
memory[15846]=8'b11111111;
memory[15847]=8'b11111111;
memory[15848]=8'b11111111;
memory[15849]=8'b11111111;
memory[15850]=8'b11111111;
memory[15851]=8'b11111111;
memory[15852]=8'b11111111;
memory[15853]=8'b11111111;
memory[15854]=8'b11111111;
memory[15855]=8'b11111111;
memory[15856]=8'b11111111;
memory[15857]=8'b11111111;
memory[15858]=8'b11111111;
memory[15859]=8'b11111111;
memory[15860]=8'b11111111;
memory[15861]=8'b11111111;
memory[15862]=8'b11111111;
memory[15863]=8'b11111111;
memory[15864]=8'b11111111;
memory[15865]=8'b11111111;
memory[15866]=8'b11111111;
memory[15867]=8'b11111111;
memory[15868]=8'b11111111;
memory[15869]=8'b11111111;
memory[15870]=8'b11111111;
memory[15871]=8'b11111111;
memory[15872]=8'b11111111;
memory[15873]=8'b11111111;
memory[15874]=8'b11111111;
memory[15875]=8'b11111111;
memory[15876]=8'b11111111;
memory[15877]=8'b11111111;
memory[15878]=8'b11111111;
memory[15879]=8'b11111111;
memory[15880]=8'b11111111;
memory[15881]=8'b11111111;
memory[15882]=8'b11111111;
memory[15883]=8'b11111111;
memory[15884]=8'b11111111;
memory[15885]=8'b11111111;
memory[15886]=8'b11111111;
memory[15887]=8'b11111111;
memory[15888]=8'b11111111;
memory[15889]=8'b11111111;
memory[15890]=8'b11111111;
memory[15891]=8'b11111111;
memory[15892]=8'b11111111;
memory[15893]=8'b11111111;
memory[15894]=8'b11111111;
memory[15895]=8'b11111111;
memory[15896]=8'b11111111;
memory[15897]=8'b11111111;
memory[15898]=8'b11111111;
memory[15899]=8'b11111111;
memory[15900]=8'b11111111;
memory[15901]=8'b11111111;
memory[15902]=8'b11111111;
memory[15903]=8'b11111111;
memory[15904]=8'b11111111;
memory[15905]=8'b11111111;
memory[15906]=8'b11111111;
memory[15907]=8'b11111111;
memory[15908]=8'b11111111;
memory[15909]=8'b11111111;
memory[15910]=8'b11111111;
memory[15911]=8'b11111111;
memory[15912]=8'b11111111;
memory[15913]=8'b11111111;
memory[15914]=8'b11111111;
memory[15915]=8'b11111111;
memory[15916]=8'b11111111;
memory[15917]=8'b11111111;
memory[15918]=8'b11111111;
memory[15919]=8'b11111111;
memory[15920]=8'b11111111;
memory[15921]=8'b11111111;
memory[15922]=8'b11111111;
memory[15923]=8'b11111111;
memory[15924]=8'b11111111;
memory[15925]=8'b11111111;
memory[15926]=8'b11111111;
memory[15927]=8'b11111111;
memory[15928]=8'b11111111;
memory[15929]=8'b11111111;
memory[15930]=8'b11111111;
memory[15931]=8'b11111111;
memory[15932]=8'b11111111;
memory[15933]=8'b11111111;
memory[15934]=8'b11111111;
memory[15935]=8'b11111111;
memory[15936]=8'b11111111;
memory[15937]=8'b11111111;
memory[15938]=8'b11111111;
memory[15939]=8'b11111111;
memory[15940]=8'b11111111;
memory[15941]=8'b11111111;
memory[15942]=8'b11111111;
memory[15943]=8'b11111111;
memory[15944]=8'b11111111;
memory[15945]=8'b11111111;
memory[15946]=8'b11111111;
memory[15947]=8'b11111111;
memory[15948]=8'b11111111;
memory[15949]=8'b11111111;
memory[15950]=8'b11111111;
memory[15951]=8'b11111111;
memory[15952]=8'b11111111;
memory[15953]=8'b11111111;
memory[15954]=8'b11111111;
memory[15955]=8'b11111111;
memory[15956]=8'b11111111;
memory[15957]=8'b11111111;
memory[15958]=8'b11111111;
memory[15959]=8'b11111111;
memory[15960]=8'b11111111;
memory[15961]=8'b11111111;
memory[15962]=8'b11111111;
memory[15963]=8'b11111111;
memory[15964]=8'b11111111;
memory[15965]=8'b11111111;
memory[15966]=8'b11111111;
memory[15967]=8'b11111111;
memory[15968]=8'b11111111;
memory[15969]=8'b11111111;
memory[15970]=8'b11111111;
memory[15971]=8'b11111111;
memory[15972]=8'b11111111;
memory[15973]=8'b11111111;
memory[15974]=8'b11111111;
memory[15975]=8'b11111111;
memory[15976]=8'b11111111;
memory[15977]=8'b11111111;
memory[15978]=8'b11111111;
memory[15979]=8'b11111111;
memory[15980]=8'b11111111;
memory[15981]=8'b11111111;
memory[15982]=8'b11111111;
memory[15983]=8'b11111111;
memory[15984]=8'b11111111;
memory[15985]=8'b11111111;
memory[15986]=8'b11111111;
memory[15987]=8'b11111111;
memory[15988]=8'b11111111;
memory[15989]=8'b11111111;
memory[15990]=8'b11111111;
memory[15991]=8'b11111111;
memory[15992]=8'b11111111;
memory[15993]=8'b11111111;
memory[15994]=8'b11111111;
memory[15995]=8'b11111111;
memory[15996]=8'b11111111;
memory[15997]=8'b11111111;
memory[15998]=8'b11111111;
memory[15999]=8'b11111111;

//*/
  end

  always @(posedge CLK) begin
    if (WE)
      memory[Address] <= DataIn;
    else
      DataOut <= memory[Address];
  end

endmodule
